magic
tech sky130B
magscale 1 2
timestamp 1761071203
<< nwell >>
rect 1066 2159 38862 697425
<< obsli1 >>
rect 1104 2159 38824 697425
<< obsm1 >>
rect 842 2128 38824 697456
<< obsm2 >>
rect 846 2139 35242 697445
<< metal3 >>
rect 0 687352 800 687472
rect 0 667496 800 667616
rect 0 647640 800 647760
rect 0 627784 800 627904
rect 0 607928 800 608048
rect 0 588072 800 588192
rect 0 568216 800 568336
rect 0 548360 800 548480
rect 0 528504 800 528624
rect 0 508648 800 508768
rect 0 488792 800 488912
rect 0 468936 800 469056
rect 0 449080 800 449200
rect 0 429224 800 429344
rect 0 409368 800 409488
rect 0 389512 800 389632
rect 0 369656 800 369776
rect 0 349800 800 349920
rect 0 329944 800 330064
rect 0 310088 800 310208
rect 0 290232 800 290352
rect 0 270376 800 270496
rect 0 250520 800 250640
rect 0 230664 800 230784
rect 0 210808 800 210928
rect 0 190952 800 191072
rect 0 171096 800 171216
rect 0 151240 800 151360
rect 0 131384 800 131504
rect 0 111528 800 111648
rect 0 91672 800 91792
rect 0 71816 800 71936
rect 0 51960 800 52080
rect 0 32104 800 32224
rect 0 12248 800 12368
<< obsm3 >>
rect 798 687552 35246 697441
rect 880 687272 35246 687552
rect 798 667696 35246 687272
rect 880 667416 35246 667696
rect 798 647840 35246 667416
rect 880 647560 35246 647840
rect 798 627984 35246 647560
rect 880 627704 35246 627984
rect 798 608128 35246 627704
rect 880 607848 35246 608128
rect 798 588272 35246 607848
rect 880 587992 35246 588272
rect 798 568416 35246 587992
rect 880 568136 35246 568416
rect 798 548560 35246 568136
rect 880 548280 35246 548560
rect 798 528704 35246 548280
rect 880 528424 35246 528704
rect 798 508848 35246 528424
rect 880 508568 35246 508848
rect 798 488992 35246 508568
rect 880 488712 35246 488992
rect 798 469136 35246 488712
rect 880 468856 35246 469136
rect 798 449280 35246 468856
rect 880 449000 35246 449280
rect 798 429424 35246 449000
rect 880 429144 35246 429424
rect 798 409568 35246 429144
rect 880 409288 35246 409568
rect 798 389712 35246 409288
rect 880 389432 35246 389712
rect 798 369856 35246 389432
rect 880 369576 35246 369856
rect 798 350000 35246 369576
rect 880 349720 35246 350000
rect 798 330144 35246 349720
rect 880 329864 35246 330144
rect 798 310288 35246 329864
rect 880 310008 35246 310288
rect 798 290432 35246 310008
rect 880 290152 35246 290432
rect 798 270576 35246 290152
rect 880 270296 35246 270576
rect 798 250720 35246 270296
rect 880 250440 35246 250720
rect 798 230864 35246 250440
rect 880 230584 35246 230864
rect 798 211008 35246 230584
rect 880 210728 35246 211008
rect 798 191152 35246 210728
rect 880 190872 35246 191152
rect 798 171296 35246 190872
rect 880 171016 35246 171296
rect 798 151440 35246 171016
rect 880 151160 35246 151440
rect 798 131584 35246 151160
rect 880 131304 35246 131584
rect 798 111728 35246 131304
rect 880 111448 35246 111728
rect 798 91872 35246 111448
rect 880 91592 35246 91872
rect 798 72016 35246 91592
rect 880 71736 35246 72016
rect 798 52160 35246 71736
rect 880 51880 35246 52160
rect 798 32304 35246 51880
rect 880 32024 35246 32304
rect 798 12448 35246 32024
rect 880 12168 35246 12448
rect 798 2143 35246 12168
<< metal4 >>
rect 4208 2128 4528 697456
rect 19568 2128 19888 697456
rect 34928 2128 35248 697456
<< obsm4 >>
rect 6499 12275 8589 323781
<< labels >>
rlabel metal3 s 0 51960 800 52080 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 647640 800 647760 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 0 171096 800 171216 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 0 230664 800 230784 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 0 290232 800 290352 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 0 349800 800 349920 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 0 409368 800 409488 6 io_in[6]
port 8 nsew signal input
rlabel metal3 s 0 468936 800 469056 6 io_in[7]
port 9 nsew signal input
rlabel metal3 s 0 528504 800 528624 6 io_in[8]
port 10 nsew signal input
rlabel metal3 s 0 588072 800 588192 6 io_in[9]
port 11 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 io_oeb[0]
port 12 nsew signal output
rlabel metal3 s 0 687352 800 687472 6 io_oeb[10]
port 13 nsew signal output
rlabel metal3 s 0 151240 800 151360 6 io_oeb[1]
port 14 nsew signal output
rlabel metal3 s 0 210808 800 210928 6 io_oeb[2]
port 15 nsew signal output
rlabel metal3 s 0 270376 800 270496 6 io_oeb[3]
port 16 nsew signal output
rlabel metal3 s 0 329944 800 330064 6 io_oeb[4]
port 17 nsew signal output
rlabel metal3 s 0 389512 800 389632 6 io_oeb[5]
port 18 nsew signal output
rlabel metal3 s 0 449080 800 449200 6 io_oeb[6]
port 19 nsew signal output
rlabel metal3 s 0 508648 800 508768 6 io_oeb[7]
port 20 nsew signal output
rlabel metal3 s 0 568216 800 568336 6 io_oeb[8]
port 21 nsew signal output
rlabel metal3 s 0 627784 800 627904 6 io_oeb[9]
port 22 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 io_out[0]
port 23 nsew signal output
rlabel metal3 s 0 667496 800 667616 6 io_out[10]
port 24 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 io_out[1]
port 25 nsew signal output
rlabel metal3 s 0 190952 800 191072 6 io_out[2]
port 26 nsew signal output
rlabel metal3 s 0 250520 800 250640 6 io_out[3]
port 27 nsew signal output
rlabel metal3 s 0 310088 800 310208 6 io_out[4]
port 28 nsew signal output
rlabel metal3 s 0 369656 800 369776 6 io_out[5]
port 29 nsew signal output
rlabel metal3 s 0 429224 800 429344 6 io_out[6]
port 30 nsew signal output
rlabel metal3 s 0 488792 800 488912 6 io_out[7]
port 31 nsew signal output
rlabel metal3 s 0 548360 800 548480 6 io_out[8]
port 32 nsew signal output
rlabel metal3 s 0 607928 800 608048 6 io_out[9]
port 33 nsew signal output
rlabel metal4 s 4208 2128 4528 697456 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 697456 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 697456 6 vssd1
port 35 nsew ground bidirectional
rlabel metal3 s 0 12248 800 12368 6 wb_clk_i
port 36 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 wb_rst_i
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 700000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9092472
string GDS_FILE /home/ghp7482/projects/LLM4Microwatt/openlane/user_proj_timer/runs/25_10_21_14_24/results/signoff/user_proj_timer.magic.gds
string GDS_START 483906
<< end >>

