magic
tech sky130B
magscale 1 2
timestamp 1761071591
<< nwell >>
rect 571138 49159 608934 744425
<< obsli1 >>
rect 571176 49159 608896 744425
<< obsm1 >>
rect 566 8 609158 953284
<< metal2 >>
rect 27498 953270 27558 953726
rect 29498 953270 29558 953726
rect 34360 953270 34416 953726
rect 34912 953270 34968 953726
rect 35556 953270 35612 953726
rect 36200 953270 36256 953726
rect 38040 953270 38096 953726
rect 38592 953270 38648 953726
rect 39236 953270 39292 953726
rect 39880 953270 39936 953726
rect 42364 953270 42420 953726
rect 42916 953270 42972 953726
rect 43560 953270 43616 953726
rect 44204 953270 44260 953726
rect 44677 953270 44891 953726
rect 45400 953270 45456 953726
rect 46560 953270 46688 953726
rect 47240 953270 47296 953726
rect 49080 953270 49136 953726
rect 78698 953270 78758 953726
rect 80698 953270 80758 953726
rect 85760 953270 85816 953726
rect 86312 953270 86368 953726
rect 86956 953270 87012 953726
rect 87600 953270 87656 953726
rect 89440 953270 89496 953726
rect 89992 953270 90048 953726
rect 90636 953270 90692 953726
rect 91280 953270 91336 953726
rect 93764 953270 93820 953726
rect 94316 953270 94372 953726
rect 94960 953270 95016 953726
rect 95604 953270 95660 953726
rect 96077 953270 96291 953726
rect 96800 953270 96856 953726
rect 97960 953270 98088 953726
rect 98640 953270 98696 953726
rect 100480 953270 100536 953726
rect 129898 953270 129958 953726
rect 131898 953270 131958 953726
rect 137160 953270 137216 953726
rect 137712 953270 137768 953726
rect 138356 953270 138412 953726
rect 139000 953270 139056 953726
rect 140840 953270 140896 953726
rect 141392 953270 141448 953726
rect 142036 953270 142092 953726
rect 142680 953270 142736 953726
rect 145164 953270 145220 953726
rect 145716 953244 145772 953726
rect 146360 953270 146416 953726
rect 147004 953270 147060 953726
rect 147477 953270 147691 953726
rect 148200 953270 148256 953726
rect 149360 953270 149488 953726
rect 150040 953270 150096 953726
rect 151880 953270 151936 953726
rect 181098 953270 181158 953726
rect 183098 953270 183158 953726
rect 188560 953270 188616 953726
rect 189112 953270 189168 953726
rect 189756 953270 189812 953726
rect 190400 953270 190456 953726
rect 192240 953270 192296 953726
rect 192792 953270 192848 953726
rect 193436 953270 193492 953726
rect 194080 953270 194136 953726
rect 196564 953270 196620 953726
rect 197116 953270 197172 953726
rect 197760 953270 197816 953726
rect 198404 953270 198460 953726
rect 198877 953270 199091 953726
rect 199600 953270 199656 953726
rect 200760 953270 200888 953726
rect 201440 953270 201496 953726
rect 203280 953270 203336 953726
rect 232298 953270 232358 953726
rect 234298 953270 234358 953726
rect 240160 953270 240216 953726
rect 240712 953270 240768 953726
rect 241356 953270 241412 953726
rect 242000 953270 242056 953726
rect 243840 953270 243896 953726
rect 244392 953244 244448 953726
rect 245036 953270 245092 953726
rect 245680 953244 245736 953726
rect 248164 953270 248220 953726
rect 248716 953270 248772 953726
rect 249360 953270 249416 953726
rect 250004 953270 250060 953726
rect 250477 953270 250691 953726
rect 251200 953270 251256 953726
rect 252360 953270 252488 953726
rect 253040 953270 253096 953726
rect 254880 953270 254936 953726
rect 336698 953270 336758 953726
rect 338698 953270 338758 953726
rect 341960 953270 342016 953726
rect 342512 953270 342568 953726
rect 343156 953270 343212 953726
rect 343800 953270 343856 953726
rect 345640 953270 345696 953726
rect 346192 953270 346248 953726
rect 346836 953270 346892 953726
rect 347480 953270 347536 953726
rect 349964 953270 350020 953726
rect 350516 953270 350572 953726
rect 351160 953270 351216 953726
rect 351804 953270 351860 953726
rect 352277 953270 352491 953726
rect 353000 953270 353056 953726
rect 354160 953270 354288 953726
rect 354840 953270 354896 953726
rect 356680 953270 356736 953726
rect 425698 953270 425758 953726
rect 427698 953270 427758 953726
rect 430960 953270 431016 953726
rect 431512 953270 431568 953726
rect 432156 953270 432212 953726
rect 432800 953270 432856 953726
rect 434640 953270 434696 953726
rect 435192 953270 435248 953726
rect 435836 953270 435892 953726
rect 436480 953270 436536 953726
rect 438964 953270 439020 953726
rect 439516 953270 439572 953726
rect 440160 953270 440216 953726
rect 440804 953270 440860 953726
rect 441277 953270 441491 953726
rect 442000 953270 442056 953726
rect 443160 953270 443288 953726
rect 443840 953270 443896 953726
rect 445680 953270 445736 953726
rect 476898 953270 476958 953726
rect 478898 953270 478958 953726
rect 482360 953270 482416 953726
rect 482912 953270 482968 953726
rect 483556 953270 483612 953726
rect 484200 953270 484256 953726
rect 486040 953270 486096 953726
rect 486592 953270 486648 953726
rect 487236 953270 487292 953726
rect 487880 953270 487936 953726
rect 490364 953270 490420 953726
rect 490916 953270 490972 953726
rect 491560 953270 491616 953726
rect 492204 953270 492260 953726
rect 492677 953270 492891 953726
rect 493400 953270 493456 953726
rect 494560 953270 494688 953726
rect 495240 953270 495296 953726
rect 497080 953270 497136 953726
rect 576298 953270 576358 953726
rect 578298 953270 578358 953726
rect 584160 953270 584216 953726
rect 584712 953270 584768 953726
rect 585356 953270 585412 953726
rect 586000 953270 586056 953726
rect 587840 953270 587896 953726
rect 588392 953270 588448 953726
rect 589036 953270 589092 953726
rect 589680 953270 589736 953726
rect 592164 953270 592220 953726
rect 592716 953270 592772 953726
rect 593360 953270 593416 953726
rect 594004 953270 594060 953726
rect 594477 953270 594691 953726
rect 595200 953270 595256 953726
rect 596360 953270 596488 953726
rect 597040 953270 597096 953726
rect 598880 953270 598936 953726
rect 99576 -400 99632 56
rect 110164 -400 110220 56
rect 145190 -400 145246 56
rect 147030 -400 147086 56
rect 147638 -400 147766 56
rect 148870 -400 148926 56
rect 149435 -400 149649 56
rect 150066 -400 150122 56
rect 150710 -400 150766 56
rect 151354 -400 151410 56
rect 151906 -400 151962 56
rect 154390 -400 154446 56
rect 155034 -400 155090 56
rect 155678 -400 155734 56
rect 156230 -400 156286 56
rect 158070 -400 158126 56
rect 158714 -400 158770 56
rect 159358 -400 159414 56
rect 159910 -400 159966 56
rect 160580 -400 160632 56
rect 163791 -400 163843 56
rect 253790 -400 253846 56
rect 255630 -400 255686 56
rect 256238 -400 256366 56
rect 257470 -400 257526 56
rect 258035 -400 258249 56
rect 258666 -400 258722 56
rect 259310 -400 259366 56
rect 259954 -400 260010 56
rect 260506 -400 260562 56
rect 262990 -400 263046 56
rect 263634 -400 263690 56
rect 264278 -400 264334 56
rect 264830 -400 264886 56
rect 266670 -400 266726 56
rect 267314 -400 267370 56
rect 267958 -400 268014 56
rect 268510 -400 268566 56
rect 269180 -400 269232 56
rect 273360 -400 273412 56
rect 308590 -400 308646 56
rect 310430 -400 310486 56
rect 311038 -400 311166 56
rect 312270 -400 312326 56
rect 312835 -400 313049 56
rect 313466 -400 313522 56
rect 314110 -400 314166 56
rect 314754 -400 314810 56
rect 315306 -400 315362 56
rect 317790 -400 317846 56
rect 318434 -400 318490 56
rect 319078 -400 319134 56
rect 319630 -400 319686 56
rect 321470 -400 321526 56
rect 322114 -400 322170 56
rect 322758 -400 322814 56
rect 323310 -400 323366 56
rect 323980 -400 324032 56
rect 328165 -400 328217 56
rect 363390 -400 363446 56
rect 365230 -400 365286 56
rect 365838 -400 365966 56
rect 367070 -400 367126 56
rect 367635 -400 367849 56
rect 368266 -400 368322 56
rect 368910 -400 368966 56
rect 369554 -400 369610 56
rect 370106 -400 370162 56
rect 372590 -400 372646 56
rect 373234 -400 373290 56
rect 373878 -400 373934 56
rect 374430 -400 374486 56
rect 376270 -400 376326 56
rect 376914 -400 376970 56
rect 377558 -400 377614 56
rect 378110 -400 378166 56
rect 378780 -400 378832 56
rect 382978 -400 383030 56
rect 418190 -400 418246 56
rect 420030 -400 420086 56
rect 420638 -400 420766 56
rect 421870 -400 421926 56
rect 422435 -400 422649 56
rect 423066 -400 423122 56
rect 423710 -400 423766 56
rect 424354 -400 424410 56
rect 424906 -400 424962 56
rect 427390 -400 427446 56
rect 428034 -400 428090 56
rect 428678 -400 428734 56
rect 429230 -400 429286 56
rect 431070 -400 431126 56
rect 431714 -400 431770 56
rect 432358 -400 432414 56
rect 432910 -400 432966 56
rect 433580 -400 433632 56
rect 437778 -400 437830 56
rect 472990 -400 473046 56
rect 474830 -400 474886 56
rect 475438 -400 475566 56
rect 476670 -400 476726 56
rect 477235 -400 477449 56
rect 477866 -400 477922 56
rect 478510 -400 478566 56
rect 479154 -400 479210 56
rect 479706 -400 479762 56
rect 482190 -400 482246 56
rect 482834 -400 482890 56
rect 483478 -400 483534 56
rect 484030 -400 484086 56
rect 485870 -400 485926 56
rect 486514 -400 486570 56
rect 487158 -400 487214 56
rect 487710 -400 487766 56
rect 488380 -400 488432 56
rect 492635 -400 492687 56
rect 605082 -400 605134 56
rect 605306 -400 605358 56
rect 605530 -400 605582 56
rect 605754 -400 605806 56
rect 605978 -400 606030 56
rect 606202 -400 606254 56
rect 606426 -400 606478 56
rect 606650 -400 606702 56
rect 606874 -400 606926 56
rect 607098 -400 607150 56
rect 607322 -400 607374 56
rect 607546 -400 607598 56
rect 607770 -400 607822 56
rect 607994 -400 608046 56
rect 608218 -400 608270 56
rect 608442 -400 608494 56
rect 608666 -400 608718 56
rect 608890 -400 608942 56
rect 609114 -400 609166 56
rect 609338 -400 609390 56
rect 609562 -400 609614 56
rect 609786 -400 609838 56
rect 610010 -400 610062 56
rect 610234 -400 610286 56
rect 610458 -400 610510 56
rect 610682 -400 610734 56
rect 610906 -400 610958 56
rect 611130 -400 611182 56
rect 611354 -400 611406 56
rect 611578 -400 611630 56
rect 611802 -400 611854 56
rect 612026 -400 612078 56
<< obsm2 >>
rect 18 953214 27442 953306
rect 27614 953214 29442 953306
rect 29614 953214 34304 953306
rect 34472 953214 34856 953306
rect 35024 953214 35500 953306
rect 35668 953214 36144 953306
rect 36312 953214 37984 953306
rect 38152 953214 38536 953306
rect 38704 953214 39180 953306
rect 39348 953214 39824 953306
rect 39992 953214 42308 953306
rect 42476 953214 42860 953306
rect 43028 953214 43504 953306
rect 43672 953214 44148 953306
rect 44316 953214 44621 953306
rect 44947 953214 45344 953306
rect 45512 953214 46504 953306
rect 46744 953214 47184 953306
rect 47352 953214 49024 953306
rect 49192 953214 78642 953306
rect 78814 953214 80642 953306
rect 80814 953214 85704 953306
rect 85872 953214 86256 953306
rect 86424 953214 86900 953306
rect 87068 953214 87544 953306
rect 87712 953214 89384 953306
rect 89552 953214 89936 953306
rect 90104 953214 90580 953306
rect 90748 953214 91224 953306
rect 91392 953214 93708 953306
rect 93876 953214 94260 953306
rect 94428 953214 94904 953306
rect 95072 953214 95548 953306
rect 95716 953214 96021 953306
rect 96347 953214 96744 953306
rect 96912 953214 97904 953306
rect 98144 953214 98584 953306
rect 98752 953214 100424 953306
rect 100592 953214 129842 953306
rect 130014 953214 131842 953306
rect 132014 953214 137104 953306
rect 137272 953214 137656 953306
rect 137824 953214 138300 953306
rect 138468 953214 138944 953306
rect 139112 953214 140784 953306
rect 140952 953214 141336 953306
rect 141504 953214 141980 953306
rect 142148 953214 142624 953306
rect 142792 953214 145108 953306
rect 145276 953214 145660 953306
rect 18 953188 145660 953214
rect 145828 953214 146304 953306
rect 146472 953214 146948 953306
rect 147116 953214 147421 953306
rect 147747 953214 148144 953306
rect 148312 953214 149304 953306
rect 149544 953214 149984 953306
rect 150152 953214 151824 953306
rect 151992 953214 181042 953306
rect 181214 953214 183042 953306
rect 183214 953214 188504 953306
rect 188672 953214 189056 953306
rect 189224 953214 189700 953306
rect 189868 953214 190344 953306
rect 190512 953214 192184 953306
rect 192352 953214 192736 953306
rect 192904 953214 193380 953306
rect 193548 953214 194024 953306
rect 194192 953214 196508 953306
rect 196676 953214 197060 953306
rect 197228 953214 197704 953306
rect 197872 953214 198348 953306
rect 198516 953214 198821 953306
rect 199147 953214 199544 953306
rect 199712 953214 200704 953306
rect 200944 953214 201384 953306
rect 201552 953214 203224 953306
rect 203392 953214 232242 953306
rect 232414 953214 234242 953306
rect 234414 953214 240104 953306
rect 240272 953214 240656 953306
rect 240824 953214 241300 953306
rect 241468 953214 241944 953306
rect 242112 953214 243784 953306
rect 243952 953214 244336 953306
rect 145828 953188 244336 953214
rect 244504 953214 244980 953306
rect 245148 953214 245624 953306
rect 244504 953188 245624 953214
rect 245792 953214 248108 953306
rect 248276 953214 248660 953306
rect 248828 953214 249304 953306
rect 249472 953214 249948 953306
rect 250116 953214 250421 953306
rect 250747 953214 251144 953306
rect 251312 953214 252304 953306
rect 252544 953214 252984 953306
rect 253152 953214 254824 953306
rect 254992 953214 336642 953306
rect 336814 953214 338642 953306
rect 338814 953214 341904 953306
rect 342072 953214 342456 953306
rect 342624 953214 343100 953306
rect 343268 953214 343744 953306
rect 343912 953214 345584 953306
rect 345752 953214 346136 953306
rect 346304 953214 346780 953306
rect 346948 953214 347424 953306
rect 347592 953214 349908 953306
rect 350076 953214 350460 953306
rect 350628 953214 351104 953306
rect 351272 953214 351748 953306
rect 351916 953214 352221 953306
rect 352547 953214 352944 953306
rect 353112 953214 354104 953306
rect 354344 953214 354784 953306
rect 354952 953214 356624 953306
rect 356792 953214 425642 953306
rect 425814 953214 427642 953306
rect 427814 953214 430904 953306
rect 431072 953214 431456 953306
rect 431624 953214 432100 953306
rect 432268 953214 432744 953306
rect 432912 953214 434584 953306
rect 434752 953214 435136 953306
rect 435304 953214 435780 953306
rect 435948 953214 436424 953306
rect 436592 953214 438908 953306
rect 439076 953214 439460 953306
rect 439628 953214 440104 953306
rect 440272 953214 440748 953306
rect 440916 953214 441221 953306
rect 441547 953214 441944 953306
rect 442112 953214 443104 953306
rect 443344 953214 443784 953306
rect 443952 953214 445624 953306
rect 445792 953214 476842 953306
rect 477014 953214 478842 953306
rect 479014 953214 482304 953306
rect 482472 953214 482856 953306
rect 483024 953214 483500 953306
rect 483668 953214 484144 953306
rect 484312 953214 485984 953306
rect 486152 953214 486536 953306
rect 486704 953214 487180 953306
rect 487348 953214 487824 953306
rect 487992 953214 490308 953306
rect 490476 953214 490860 953306
rect 491028 953214 491504 953306
rect 491672 953214 492148 953306
rect 492316 953214 492621 953306
rect 492947 953214 493344 953306
rect 493512 953214 494504 953306
rect 494744 953214 495184 953306
rect 495352 953214 497024 953306
rect 497192 953214 576242 953306
rect 576414 953214 578242 953306
rect 578414 953214 584104 953306
rect 584272 953214 584656 953306
rect 584824 953214 585300 953306
rect 585468 953214 585944 953306
rect 586112 953214 587784 953306
rect 587952 953214 588336 953306
rect 588504 953214 588980 953306
rect 589148 953214 589624 953306
rect 589792 953214 592108 953306
rect 592276 953214 592660 953306
rect 592828 953214 593304 953306
rect 593472 953214 593948 953306
rect 594116 953214 594421 953306
rect 594747 953214 595144 953306
rect 595312 953214 596304 953306
rect 596544 953214 596984 953306
rect 597152 953214 598824 953306
rect 598992 953214 633310 953306
rect 245792 953188 633310 953214
rect 18 112 633310 953188
rect 18 2 99520 112
rect 99688 2 110108 112
rect 110276 2 145134 112
rect 145302 2 146974 112
rect 147142 2 147582 112
rect 147822 2 148814 112
rect 148982 2 149379 112
rect 149705 2 150010 112
rect 150178 2 150654 112
rect 150822 2 151298 112
rect 151466 2 151850 112
rect 152018 2 154334 112
rect 154502 2 154978 112
rect 155146 2 155622 112
rect 155790 2 156174 112
rect 156342 2 158014 112
rect 158182 2 158658 112
rect 158826 2 159302 112
rect 159470 2 159854 112
rect 160022 2 160524 112
rect 160688 2 163735 112
rect 163899 2 253734 112
rect 253902 2 255574 112
rect 255742 2 256182 112
rect 256422 2 257414 112
rect 257582 2 257979 112
rect 258305 2 258610 112
rect 258778 2 259254 112
rect 259422 2 259898 112
rect 260066 2 260450 112
rect 260618 2 262934 112
rect 263102 2 263578 112
rect 263746 2 264222 112
rect 264390 2 264774 112
rect 264942 2 266614 112
rect 266782 2 267258 112
rect 267426 2 267902 112
rect 268070 2 268454 112
rect 268622 2 269124 112
rect 269288 2 273304 112
rect 273468 2 308534 112
rect 308702 2 310374 112
rect 310542 2 310982 112
rect 311222 2 312214 112
rect 312382 2 312779 112
rect 313105 2 313410 112
rect 313578 2 314054 112
rect 314222 2 314698 112
rect 314866 2 315250 112
rect 315418 2 317734 112
rect 317902 2 318378 112
rect 318546 2 319022 112
rect 319190 2 319574 112
rect 319742 2 321414 112
rect 321582 2 322058 112
rect 322226 2 322702 112
rect 322870 2 323254 112
rect 323422 2 323924 112
rect 324088 2 328109 112
rect 328273 2 363334 112
rect 363502 2 365174 112
rect 365342 2 365782 112
rect 366022 2 367014 112
rect 367182 2 367579 112
rect 367905 2 368210 112
rect 368378 2 368854 112
rect 369022 2 369498 112
rect 369666 2 370050 112
rect 370218 2 372534 112
rect 372702 2 373178 112
rect 373346 2 373822 112
rect 373990 2 374374 112
rect 374542 2 376214 112
rect 376382 2 376858 112
rect 377026 2 377502 112
rect 377670 2 378054 112
rect 378222 2 378724 112
rect 378888 2 382922 112
rect 383086 2 418134 112
rect 418302 2 419974 112
rect 420142 2 420582 112
rect 420822 2 421814 112
rect 421982 2 422379 112
rect 422705 2 423010 112
rect 423178 2 423654 112
rect 423822 2 424298 112
rect 424466 2 424850 112
rect 425018 2 427334 112
rect 427502 2 427978 112
rect 428146 2 428622 112
rect 428790 2 429174 112
rect 429342 2 431014 112
rect 431182 2 431658 112
rect 431826 2 432302 112
rect 432470 2 432854 112
rect 433022 2 433524 112
rect 433688 2 437722 112
rect 437886 2 472934 112
rect 473102 2 474774 112
rect 474942 2 475382 112
rect 475622 2 476614 112
rect 476782 2 477179 112
rect 477505 2 477810 112
rect 477978 2 478454 112
rect 478622 2 479098 112
rect 479266 2 479650 112
rect 479818 2 482134 112
rect 482302 2 482778 112
rect 482946 2 483422 112
rect 483590 2 483974 112
rect 484142 2 485814 112
rect 485982 2 486458 112
rect 486626 2 487102 112
rect 487270 2 487654 112
rect 487822 2 488324 112
rect 488488 2 492579 112
rect 492743 2 605026 112
rect 605190 2 605250 112
rect 605414 2 605474 112
rect 605638 2 605698 112
rect 605862 2 605922 112
rect 606086 2 606146 112
rect 606310 2 606370 112
rect 606534 2 606594 112
rect 606758 2 606818 112
rect 606982 2 607042 112
rect 607206 2 607266 112
rect 607430 2 607490 112
rect 607654 2 607714 112
rect 607878 2 607938 112
rect 608102 2 608162 112
rect 608326 2 608386 112
rect 608550 2 608610 112
rect 608774 2 608834 112
rect 608998 2 609058 112
rect 609222 2 609282 112
rect 609446 2 609506 112
rect 609670 2 609730 112
rect 609894 2 609954 112
rect 610118 2 610178 112
rect 610342 2 610402 112
rect 610566 2 610626 112
rect 610790 2 610850 112
rect 611014 2 611074 112
rect 611238 2 611298 112
rect 611462 2 611522 112
rect 611686 2 611746 112
rect 611910 2 611970 112
rect 612134 2 633310 112
<< metal3 >>
rect 291362 953266 296142 953726
rect 301342 953266 306122 953726
rect 533562 953266 538342 953726
rect 543542 953266 548322 953726
rect 633266 929006 633726 929068
rect -400 927072 60 927142
rect 633266 927006 633726 927068
rect -400 925232 60 925302
rect 633266 925104 633726 925174
rect -400 924560 60 924688
rect 633266 924552 633726 924622
rect 633266 923908 633726 923978
rect -400 923392 60 923462
rect 633266 923264 633726 923334
rect -400 922677 60 922891
rect -400 922196 60 922266
rect -400 921552 60 921622
rect 633266 921424 633726 921494
rect -400 920908 60 920978
rect 633266 920872 633726 920942
rect -400 920356 60 920426
rect 633266 920228 633726 920298
rect 633266 919584 633726 919654
rect -400 917872 60 917942
rect -400 917228 60 917298
rect 633266 917100 633726 917170
rect -400 916584 60 916654
rect 633266 916548 633726 916618
rect -400 916032 60 916102
rect 633266 915904 633726 915974
rect 633266 915260 633726 915330
rect 633266 914635 633726 914849
rect -400 914192 60 914262
rect 633266 914064 633726 914134
rect -400 913548 60 913618
rect -400 912904 60 912974
rect 633266 912838 633726 912966
rect -400 912352 60 912422
rect 633266 912224 633726 912294
rect 633266 910384 633726 910454
rect -400 906644 60 906704
rect -400 904644 122 904704
rect -400 880014 60 884804
rect -400 875054 60 879716
rect 633571 875562 633726 880362
rect -400 869964 60 874764
rect 633571 870610 633726 875272
rect 633571 865522 633726 870312
rect -400 837742 60 842522
rect 633266 839006 633726 839068
rect 633266 837006 633726 837068
rect 633266 835904 633726 835974
rect 633266 835352 633726 835422
rect 633266 834708 633726 834778
rect 633266 834064 633726 834134
rect -400 827762 60 832542
rect 633266 832224 633726 832294
rect 633206 831672 633726 831742
rect 633266 831028 633726 831098
rect 633266 830384 633726 830454
rect 633266 827900 633726 827970
rect 633266 827348 633726 827418
rect 633266 826704 633726 826774
rect 633266 826060 633726 826130
rect 633266 825435 633726 825649
rect 633266 824864 633726 824934
rect 633266 823638 633726 823766
rect 633266 823024 633726 823094
rect 633266 821184 633726 821254
rect -400 795542 60 800322
rect -400 785562 60 790342
rect 633266 786384 633726 791164
rect 633266 776406 633726 781186
rect -400 757272 60 757342
rect -400 755432 60 755502
rect -400 754760 60 754888
rect -400 753592 60 753662
rect -400 752877 60 753091
rect -400 752396 60 752466
rect -400 751752 60 751822
rect -400 751108 60 751178
rect -400 750556 60 750626
rect 633266 750006 633726 750068
rect -400 748072 60 748142
rect 633266 748006 633726 748068
rect -400 747428 60 747498
rect -400 746784 60 746854
rect 633266 746704 633726 746774
rect -400 746232 60 746302
rect 633266 746152 633726 746222
rect 633266 745508 633726 745578
rect 633266 744864 633726 744934
rect -400 744392 60 744462
rect -400 743748 60 743818
rect -400 743104 60 743174
rect 633266 743024 633726 743094
rect -400 742552 60 742622
rect 633266 742472 633726 742542
rect 633266 741828 633726 741898
rect 633206 741184 633726 741254
rect 633266 738700 633726 738770
rect 633266 738148 633726 738218
rect 633266 737504 633726 737574
rect 633266 736860 633726 736930
rect -400 736644 60 736704
rect 633266 736235 633726 736449
rect 633266 735664 633726 735734
rect -400 734644 122 734704
rect 633266 734438 633726 734566
rect 633266 733824 633726 733894
rect 633266 731984 633726 732054
rect -400 714072 60 714142
rect -400 712232 60 712302
rect -400 711560 60 711688
rect -400 710392 60 710462
rect -400 709677 60 709891
rect -400 709196 60 709266
rect -400 708552 60 708622
rect -400 707908 60 707978
rect -400 707356 60 707426
rect -400 704872 60 704942
rect 633266 705006 633726 705068
rect -400 704228 60 704298
rect -400 703584 60 703654
rect -400 703032 60 703102
rect 633266 703006 633726 703068
rect 633266 701704 633726 701774
rect -400 701192 60 701262
rect 633266 701152 633726 701222
rect -400 700548 60 700618
rect 633266 700508 633726 700578
rect -400 699904 60 699974
rect 633266 699864 633726 699934
rect -400 699352 60 699422
rect 633266 698024 633726 698094
rect 633266 697472 633726 697542
rect 633266 696828 633726 696898
rect 633266 696184 633726 696254
rect -400 693644 60 693704
rect 633266 693700 633726 693770
rect 633266 693148 633726 693218
rect 633266 692504 633726 692574
rect 633266 691860 633726 691930
rect -400 691644 674 691704
rect 633266 691235 633726 691449
rect 633266 690664 633726 690734
rect 633266 689438 633726 689566
rect 633266 688824 633726 688894
rect 633266 686984 633726 687054
rect -400 670872 60 670942
rect -400 669032 60 669102
rect -400 668360 60 668488
rect -400 667192 60 667262
rect -400 666477 60 666691
rect -400 665996 60 666066
rect -400 665352 60 665422
rect -400 664708 60 664778
rect -400 664156 60 664226
rect -400 661672 60 661742
rect -400 661028 60 661098
rect -400 660384 60 660454
rect 633266 660006 633726 660068
rect -400 659832 60 659902
rect -400 657992 60 658062
rect 633266 658006 633726 658068
rect -400 657348 60 657418
rect -400 656704 60 656774
rect 633266 656704 633726 656774
rect -400 656152 60 656222
rect 633266 656152 633726 656222
rect 633266 655508 633726 655578
rect 633266 654864 633726 654934
rect 633266 653024 633726 653094
rect 633266 652472 633726 652542
rect 633266 651828 633726 651898
rect 633266 651184 633726 651254
rect -400 650644 60 650704
rect -400 648644 674 648704
rect 633266 648700 633726 648770
rect 633266 648148 633726 648218
rect 633266 647504 633726 647574
rect 633266 646860 633726 646930
rect 633266 646235 633726 646449
rect 633266 645664 633726 645734
rect 633266 644438 633726 644566
rect 633266 643824 633726 643894
rect 633266 641984 633726 642054
rect -400 627672 60 627742
rect -400 625832 60 625902
rect -400 625160 60 625288
rect -400 623992 60 624062
rect -400 623277 60 623491
rect -400 622796 60 622866
rect -400 622152 60 622222
rect -400 621508 60 621578
rect -400 620956 60 621026
rect -400 618472 60 618542
rect -400 617828 60 617898
rect -400 617184 60 617254
rect -400 616632 60 616702
rect 633266 615006 633726 615068
rect -400 614792 60 614862
rect -400 614148 60 614218
rect -400 613504 60 613574
rect -400 612952 60 613022
rect 633266 613006 633726 613068
rect 633266 611504 633726 611574
rect 633266 610952 633726 611022
rect 633266 610308 633726 610378
rect 633266 609664 633726 609734
rect 633266 607824 633726 607894
rect -400 607644 60 607704
rect 633266 607272 633726 607342
rect 633266 606628 633726 606698
rect 633266 605984 633726 606054
rect -400 605644 674 605704
rect 633266 603500 633726 603570
rect 633266 602948 633726 603018
rect 633266 602304 633726 602374
rect 633266 601660 633726 601730
rect 633266 601035 633726 601249
rect 633266 600464 633726 600534
rect 633266 599238 633726 599366
rect 633266 598624 633726 598694
rect 633266 596784 633726 596854
rect -400 584472 60 584542
rect -400 582632 60 582702
rect -400 581960 60 582088
rect -400 580792 60 580862
rect -400 580077 60 580291
rect -400 579596 60 579666
rect -400 578952 60 579022
rect -400 578308 60 578378
rect -400 577756 60 577826
rect -400 575272 60 575342
rect -400 574628 60 574698
rect -400 573984 60 574054
rect -400 573432 60 573502
rect -400 571592 60 571662
rect -400 570948 60 571018
rect -400 570304 60 570374
rect 633266 570006 633726 570068
rect -400 569752 60 569822
rect 633266 568006 633726 568068
rect 633266 566504 633726 566574
rect 633266 565952 633726 566022
rect 633266 565308 633726 565378
rect -400 564644 60 564704
rect 633266 564664 633726 564734
rect 633266 562824 633726 562894
rect -400 562644 674 562704
rect 633266 562272 633726 562342
rect 633266 561628 633726 561698
rect 633266 560984 633726 561054
rect 633266 558500 633726 558570
rect 633266 557948 633726 558018
rect 633266 557304 633726 557374
rect 633266 556660 633726 556730
rect 633266 556035 633726 556249
rect 633266 555464 633726 555534
rect 633266 554238 633726 554366
rect 633266 553624 633726 553694
rect 633266 551784 633726 551854
rect -400 541272 60 541342
rect -400 539432 60 539502
rect -400 538760 60 538888
rect -400 537592 60 537662
rect -400 536877 60 537091
rect -400 536396 60 536466
rect -400 535752 60 535822
rect -400 535108 60 535178
rect -400 534556 60 534626
rect -400 532072 60 532142
rect -400 531428 60 531498
rect -400 530784 60 530854
rect -400 530232 60 530302
rect -400 528392 60 528462
rect -400 527748 60 527818
rect -400 527104 60 527174
rect -400 526552 60 526622
rect 633266 525006 633726 525068
rect 633266 523005 633726 523067
rect -400 521644 60 521704
rect 633266 521304 633726 521374
rect 633266 520752 633726 520822
rect 633266 520108 633726 520178
rect -400 519644 674 519704
rect 633266 519464 633726 519534
rect 633266 517624 633726 517694
rect 633266 517072 633726 517142
rect 633266 516428 633726 516498
rect 633266 515784 633726 515854
rect 633266 513300 633726 513370
rect 633206 512748 633726 512818
rect 633266 512104 633726 512174
rect 633266 511460 633726 511530
rect 633266 510835 633726 511049
rect 633266 510264 633726 510334
rect 633266 509038 633726 509166
rect 633266 508424 633726 508494
rect 633266 506584 633726 506654
rect -400 498072 60 498142
rect -400 496232 60 496302
rect -400 495560 60 495688
rect -400 494392 60 494462
rect -400 493677 60 493891
rect -400 493196 60 493266
rect -400 492552 60 492622
rect -400 491908 60 491978
rect -400 491356 60 491426
rect -400 488872 60 488942
rect -400 488228 60 488298
rect -400 487584 60 487654
rect -400 487032 60 487102
rect -400 485192 60 485262
rect -400 484548 60 484618
rect -400 483904 60 483974
rect -400 483352 60 483422
rect -400 478644 60 478704
rect -400 476644 674 476704
rect 633266 471784 633726 476564
rect 633266 461804 633726 466584
rect -400 450940 60 455720
rect -400 440962 60 445742
rect 633571 427762 633726 432562
rect 633571 422810 633726 427472
rect 633571 417722 633726 422512
rect -400 408814 60 413604
rect -400 403862 60 408514
rect -400 398762 60 403562
rect 633266 383584 633726 388364
rect 633266 373606 633726 378386
rect -400 370472 60 370542
rect -400 368632 60 368702
rect -400 367960 60 368088
rect -400 366792 60 366862
rect -400 366077 60 366291
rect -400 365596 60 365666
rect -400 364952 60 365022
rect -400 364308 60 364378
rect -400 363756 60 363826
rect -400 361272 60 361342
rect -400 360628 60 360698
rect -400 359984 60 360054
rect -400 359432 60 359502
rect -400 357592 60 357662
rect -400 356948 60 357018
rect -400 356304 60 356374
rect -400 355752 60 355822
rect -400 349644 60 349704
rect 633266 348006 633726 348068
rect -400 347644 674 347704
rect 633266 346005 633726 346067
rect 633266 344104 633726 344174
rect 633266 343552 633726 343622
rect 633266 342908 633726 342978
rect 633266 342264 633726 342334
rect 633266 340424 633726 340494
rect 633266 339872 633726 339942
rect 633266 339228 633726 339298
rect 633266 338584 633726 338654
rect 633266 336100 633726 336170
rect 633266 335548 633726 335618
rect 633266 334904 633726 334974
rect 633266 334260 633726 334330
rect 633266 333635 633726 333849
rect 633266 333064 633726 333134
rect 633266 331838 633726 331966
rect 633266 331224 633726 331294
rect 633266 329384 633726 329454
rect -400 327272 60 327342
rect -400 325432 60 325502
rect -400 324760 60 324888
rect -400 323592 60 323662
rect -400 322877 60 323091
rect -400 322396 60 322466
rect -400 321752 60 321822
rect -400 321108 60 321178
rect -400 320556 60 320626
rect -400 318072 60 318142
rect -400 317428 60 317498
rect -400 316784 60 316854
rect -400 316232 60 316302
rect -400 314392 60 314462
rect -400 313748 60 313818
rect -400 313104 60 313174
rect -400 312552 60 312622
rect -400 306644 60 306704
rect -400 304644 674 304704
rect 633266 303006 633726 303068
rect 633266 301005 633726 301067
rect 633266 298904 633726 298974
rect 633266 298352 633726 298422
rect 633266 297708 633726 297778
rect 633266 297064 633726 297134
rect 633266 295224 633726 295294
rect 633266 294672 633726 294742
rect 633266 294028 633726 294098
rect 633206 293384 633726 293454
rect 633266 290900 633726 290970
rect 633266 290348 633726 290418
rect 633266 289704 633726 289774
rect 633266 289060 633726 289130
rect 633266 288435 633726 288649
rect 633266 287864 633726 287934
rect 633266 286638 633726 286766
rect 633266 286024 633726 286094
rect -400 284072 60 284142
rect 633266 284184 633726 284254
rect -400 282232 60 282302
rect -400 281560 60 281688
rect -400 280392 60 280462
rect -400 279677 60 279891
rect -400 279196 60 279266
rect -400 278552 60 278622
rect -400 277908 60 277978
rect -400 277356 60 277426
rect -400 274872 60 274942
rect -400 274228 60 274298
rect -400 273584 60 273654
rect -400 273032 60 273102
rect -400 271192 60 271262
rect -400 270548 60 270618
rect -400 269904 60 269974
rect -400 269352 60 269422
rect -400 263644 60 263704
rect -400 261644 674 261704
rect 633266 258006 633726 258068
rect 633266 256005 633726 256067
rect 633266 253904 633726 253974
rect 633266 253352 633726 253422
rect 633266 252708 633726 252778
rect 633266 252064 633726 252134
rect 633266 250224 633726 250294
rect 633266 249672 633726 249742
rect 633266 249028 633726 249098
rect 633266 248384 633726 248454
rect 633266 245900 633726 245970
rect 633266 245348 633726 245418
rect 633266 244704 633726 244774
rect 633266 244060 633726 244130
rect 633266 243435 633726 243649
rect 633266 242864 633726 242934
rect 633266 241638 633726 241766
rect 633266 241024 633726 241094
rect -400 240872 60 240942
rect 633266 239184 633726 239254
rect -400 239032 60 239102
rect -400 238360 60 238488
rect -400 237192 60 237262
rect -400 236477 60 236691
rect -400 235996 60 236066
rect -400 235352 60 235422
rect -400 234708 60 234778
rect -400 234156 60 234226
rect -400 231672 60 231742
rect -400 231028 60 231098
rect -400 230384 60 230454
rect -400 229832 60 229902
rect -400 227992 60 228062
rect -400 227348 60 227418
rect -400 226704 60 226774
rect -400 226152 60 226222
rect -400 220644 60 220704
rect -400 218644 674 218704
rect 633266 213006 633726 213068
rect 633266 211005 633726 211067
rect 633266 208904 633726 208974
rect 633266 208352 633726 208422
rect 633266 207708 633726 207778
rect 633266 207064 633726 207134
rect 633266 205224 633726 205294
rect 633266 204672 633726 204742
rect 633266 204028 633726 204098
rect 633266 203384 633726 203454
rect 633266 200900 633726 200970
rect 633266 200348 633726 200418
rect 633266 199704 633726 199774
rect 633266 199060 633726 199130
rect 633266 198435 633726 198649
rect 633266 197864 633726 197934
rect -400 197672 60 197742
rect 633266 196638 633726 196766
rect 633266 196024 633726 196094
rect -400 195832 60 195902
rect -400 195160 60 195288
rect 633266 194184 633726 194254
rect -400 193992 60 194062
rect -400 193277 60 193491
rect -400 192796 60 192866
rect -400 192152 60 192222
rect -400 191508 60 191578
rect -400 190956 60 191026
rect -400 188472 60 188542
rect -400 187828 60 187898
rect -400 187184 60 187254
rect -400 186632 60 186702
rect -400 184792 60 184862
rect -400 184148 60 184218
rect -400 183504 60 183574
rect -400 182952 60 183022
rect -400 177644 60 177704
rect -400 175644 674 175704
rect 633266 168006 633726 168068
rect 633266 166005 633726 166067
rect 633266 163704 633726 163774
rect 633266 163152 633726 163222
rect 633266 162508 633726 162578
rect 633266 161864 633726 161934
rect 633266 160024 633726 160094
rect 633266 159472 633726 159542
rect 633266 158828 633726 158898
rect 633266 158184 633726 158254
rect 633266 155700 633726 155770
rect 633266 155148 633726 155218
rect -400 154472 60 154542
rect 633266 154504 633726 154574
rect 633266 153860 633726 153930
rect 633266 153235 633726 153449
rect -400 152632 60 152702
rect 633266 152664 633726 152734
rect -400 151960 60 152088
rect 633266 151438 633726 151566
rect -400 150792 60 150862
rect 633266 150824 633726 150894
rect -400 150077 60 150291
rect -400 149596 60 149666
rect -400 148952 60 149022
rect 633266 148984 633726 149054
rect -400 148308 60 148378
rect -400 147756 60 147826
rect -400 145272 60 145342
rect -400 144628 60 144698
rect -400 143984 60 144054
rect -400 143432 60 143502
rect -400 141592 60 141662
rect -400 140948 60 141018
rect -400 140304 60 140374
rect -400 139752 60 139822
rect -400 134644 60 134704
rect -400 132644 674 132704
rect 633266 123006 633726 123068
rect 633266 121005 633726 121067
rect 633266 118704 633726 118774
rect 633266 118152 633726 118222
rect 633266 117508 633726 117578
rect 633266 116864 633726 116934
rect 633266 115024 633726 115094
rect 633266 114472 633726 114542
rect 633266 113828 633726 113898
rect 633266 113184 633726 113254
rect 633266 110700 633726 110770
rect 633266 110148 633726 110218
rect 633266 109504 633726 109574
rect 633266 108860 633726 108930
rect 633266 108235 633726 108449
rect 633266 107664 633726 107734
rect 633266 106438 633726 106566
rect 633266 105824 633726 105894
rect 633266 103984 633726 104054
rect -400 78140 60 82920
rect 633266 78006 633726 78068
rect 633266 76005 633726 76067
rect 633266 73504 633726 73574
rect -400 68162 60 72942
rect 633266 72952 633726 73022
rect 633266 72308 633726 72378
rect 633266 71664 633726 71734
rect 633266 69824 633726 69894
rect 633266 69272 633726 69342
rect 633266 68628 633726 68698
rect 633266 67984 633726 68054
rect 633266 65500 633726 65570
rect 633266 64948 633726 65018
rect 633266 64304 633726 64374
rect 633266 63660 633726 63730
rect 633266 63035 633726 63249
rect 633266 62464 633726 62534
rect 633266 61238 633726 61366
rect 633266 60624 633726 60694
rect 633266 58784 633726 58854
rect -400 53595 60 53665
rect -400 53372 60 53442
rect -400 53147 60 53217
rect -400 36014 60 40804
rect -400 25962 60 30762
rect 36806 -400 41586 60
rect 46784 -400 51564 60
rect 199284 -400 203914 60
rect 209164 -400 213964 60
rect 527006 -400 531786 60
rect 536984 -400 541764 60
rect 580806 -400 585586 60
rect 590784 -400 595564 60
<< obsm3 >>
rect 0 929148 633326 949381
rect 0 928926 633186 929148
rect 0 927222 633326 928926
rect 140 927148 633326 927222
rect 140 926992 633186 927148
rect 0 926926 633186 926992
rect 0 925382 633326 926926
rect 140 925254 633326 925382
rect 140 925152 633186 925254
rect 0 925024 633186 925152
rect 0 924768 633326 925024
rect 140 924702 633326 924768
rect 140 924480 633186 924702
rect 0 924472 633186 924480
rect 0 924058 633326 924472
rect 0 923828 633186 924058
rect 0 923542 633326 923828
rect 140 923414 633326 923542
rect 140 923312 633186 923414
rect 0 923184 633186 923312
rect 0 922971 633326 923184
rect 140 922597 633326 922971
rect 0 922346 633326 922597
rect 140 922116 633326 922346
rect 0 921702 633326 922116
rect 140 921574 633326 921702
rect 140 921472 633186 921574
rect 0 921344 633186 921472
rect 0 921058 633326 921344
rect 140 921022 633326 921058
rect 140 920828 633186 921022
rect 0 920792 633186 920828
rect 0 920506 633326 920792
rect 140 920378 633326 920506
rect 140 920276 633186 920378
rect 0 920148 633186 920276
rect 0 919734 633326 920148
rect 0 919504 633186 919734
rect 0 918022 633326 919504
rect 140 917792 633326 918022
rect 0 917378 633326 917792
rect 140 917250 633326 917378
rect 140 917148 633186 917250
rect 0 917020 633186 917148
rect 0 916734 633326 917020
rect 140 916698 633326 916734
rect 140 916504 633186 916698
rect 0 916468 633186 916504
rect 0 916182 633326 916468
rect 140 916054 633326 916182
rect 140 915952 633186 916054
rect 0 915824 633186 915952
rect 0 915410 633326 915824
rect 0 915180 633186 915410
rect 0 914929 633326 915180
rect 0 914555 633186 914929
rect 0 914342 633326 914555
rect 140 914214 633326 914342
rect 140 914112 633186 914214
rect 0 913984 633186 914112
rect 0 913698 633326 913984
rect 140 913468 633326 913698
rect 0 913054 633326 913468
rect 140 913046 633326 913054
rect 140 912824 633186 913046
rect 0 912758 633186 912824
rect 0 912502 633326 912758
rect 140 912374 633326 912502
rect 140 912272 633186 912374
rect 0 912144 633186 912272
rect 0 910534 633326 912144
rect 0 910304 633186 910534
rect 0 906784 633326 910304
rect 140 906564 633326 906784
rect 0 904784 633326 906564
rect 202 904564 633326 904784
rect 0 884884 633326 904564
rect 140 880442 633326 884884
rect 140 880362 633186 880442
rect 140 879934 633571 880362
rect 0 879796 633571 879934
rect 140 874974 633571 879796
rect 0 874844 633571 874974
rect 140 869884 633571 874844
rect 0 865522 633571 869884
rect 0 865442 633186 865522
rect 0 842602 633326 865442
rect 140 839148 633326 842602
rect 140 838926 633186 839148
rect 140 837662 633326 838926
rect 0 837148 633326 837662
rect 0 836926 633186 837148
rect 0 836054 633326 836926
rect 0 835824 633186 836054
rect 0 835502 633326 835824
rect 0 835272 633186 835502
rect 0 834858 633326 835272
rect 0 834628 633186 834858
rect 0 834214 633326 834628
rect 0 833984 633186 834214
rect 0 832622 633326 833984
rect 140 832374 633326 832622
rect 140 832144 633186 832374
rect 140 831822 633326 832144
rect 140 831592 633126 831822
rect 140 831178 633326 831592
rect 140 830948 633186 831178
rect 140 830534 633326 830948
rect 140 830304 633186 830534
rect 140 828050 633326 830304
rect 140 827820 633186 828050
rect 140 827682 633326 827820
rect 0 827498 633326 827682
rect 0 827268 633186 827498
rect 0 826854 633326 827268
rect 0 826624 633186 826854
rect 0 826210 633326 826624
rect 0 825980 633186 826210
rect 0 825729 633326 825980
rect 0 825355 633186 825729
rect 0 825014 633326 825355
rect 0 824784 633186 825014
rect 0 823846 633326 824784
rect 0 823558 633186 823846
rect 0 823174 633326 823558
rect 0 822944 633186 823174
rect 0 821334 633326 822944
rect 0 821104 633186 821334
rect 0 800402 633326 821104
rect 140 795462 633326 800402
rect 0 791244 633326 795462
rect 0 790422 633186 791244
rect 140 786304 633186 790422
rect 140 785482 633326 786304
rect 0 781266 633326 785482
rect 0 776326 633186 781266
rect 0 757422 633326 776326
rect 140 757192 633326 757422
rect 0 755582 633326 757192
rect 140 755352 633326 755582
rect 0 754968 633326 755352
rect 140 754680 633326 754968
rect 0 753742 633326 754680
rect 140 753512 633326 753742
rect 0 753171 633326 753512
rect 140 752797 633326 753171
rect 0 752546 633326 752797
rect 140 752316 633326 752546
rect 0 751902 633326 752316
rect 140 751672 633326 751902
rect 0 751258 633326 751672
rect 140 751028 633326 751258
rect 0 750706 633326 751028
rect 140 750476 633326 750706
rect 0 750148 633326 750476
rect 0 749926 633186 750148
rect 0 748222 633326 749926
rect 140 748148 633326 748222
rect 140 747992 633186 748148
rect 0 747926 633186 747992
rect 0 747578 633326 747926
rect 140 747348 633326 747578
rect 0 746934 633326 747348
rect 140 746854 633326 746934
rect 140 746704 633186 746854
rect 0 746624 633186 746704
rect 0 746382 633326 746624
rect 140 746302 633326 746382
rect 140 746152 633186 746302
rect 0 746072 633186 746152
rect 0 745658 633326 746072
rect 0 745428 633186 745658
rect 0 745014 633326 745428
rect 0 744784 633186 745014
rect 0 744542 633326 744784
rect 140 744312 633326 744542
rect 0 743898 633326 744312
rect 140 743668 633326 743898
rect 0 743254 633326 743668
rect 140 743174 633326 743254
rect 140 743024 633186 743174
rect 0 742944 633186 743024
rect 0 742702 633326 742944
rect 140 742622 633326 742702
rect 140 742472 633186 742622
rect 0 742392 633186 742472
rect 0 741978 633326 742392
rect 0 741748 633186 741978
rect 0 741334 633326 741748
rect 0 741104 633126 741334
rect 0 738850 633326 741104
rect 0 738620 633186 738850
rect 0 738298 633326 738620
rect 0 738068 633186 738298
rect 0 737654 633326 738068
rect 0 737424 633186 737654
rect 0 737010 633326 737424
rect 0 736784 633186 737010
rect 140 736780 633186 736784
rect 140 736564 633326 736780
rect 0 736529 633326 736564
rect 0 736155 633186 736529
rect 0 735814 633326 736155
rect 0 735584 633186 735814
rect 0 734784 633326 735584
rect 202 734646 633326 734784
rect 202 734564 633186 734646
rect 0 734358 633186 734564
rect 0 733974 633326 734358
rect 0 733744 633186 733974
rect 0 732134 633326 733744
rect 0 731904 633186 732134
rect 0 714222 633326 731904
rect 140 713992 633326 714222
rect 0 712382 633326 713992
rect 140 712152 633326 712382
rect 0 711768 633326 712152
rect 140 711480 633326 711768
rect 0 710542 633326 711480
rect 140 710312 633326 710542
rect 0 709971 633326 710312
rect 140 709597 633326 709971
rect 0 709346 633326 709597
rect 140 709116 633326 709346
rect 0 708702 633326 709116
rect 140 708472 633326 708702
rect 0 708058 633326 708472
rect 140 707828 633326 708058
rect 0 707506 633326 707828
rect 140 707276 633326 707506
rect 0 705148 633326 707276
rect 0 705022 633186 705148
rect 140 704926 633186 705022
rect 140 704792 633326 704926
rect 0 704378 633326 704792
rect 140 704148 633326 704378
rect 0 703734 633326 704148
rect 140 703504 633326 703734
rect 0 703182 633326 703504
rect 140 703148 633326 703182
rect 140 702952 633186 703148
rect 0 702926 633186 702952
rect 0 701854 633326 702926
rect 0 701624 633186 701854
rect 0 701342 633326 701624
rect 140 701302 633326 701342
rect 140 701112 633186 701302
rect 0 701072 633186 701112
rect 0 700698 633326 701072
rect 140 700658 633326 700698
rect 140 700468 633186 700658
rect 0 700428 633186 700468
rect 0 700054 633326 700428
rect 140 700014 633326 700054
rect 140 699824 633186 700014
rect 0 699784 633186 699824
rect 0 699502 633326 699784
rect 140 699272 633326 699502
rect 0 698174 633326 699272
rect 0 697944 633186 698174
rect 0 697622 633326 697944
rect 0 697392 633186 697622
rect 0 696978 633326 697392
rect 0 696748 633186 696978
rect 0 696334 633326 696748
rect 0 696104 633186 696334
rect 0 693850 633326 696104
rect 0 693784 633186 693850
rect 140 693620 633186 693784
rect 140 693564 633326 693620
rect 0 693298 633326 693564
rect 0 693068 633186 693298
rect 0 692654 633326 693068
rect 0 692424 633186 692654
rect 0 692010 633326 692424
rect 0 691784 633186 692010
rect 754 691780 633186 691784
rect 754 691564 633326 691780
rect 0 691529 633326 691564
rect 0 691155 633186 691529
rect 0 690814 633326 691155
rect 0 690584 633186 690814
rect 0 689646 633326 690584
rect 0 689358 633186 689646
rect 0 688974 633326 689358
rect 0 688744 633186 688974
rect 0 687134 633326 688744
rect 0 686904 633186 687134
rect 0 671022 633326 686904
rect 140 670792 633326 671022
rect 0 669182 633326 670792
rect 140 668952 633326 669182
rect 0 668568 633326 668952
rect 140 668280 633326 668568
rect 0 667342 633326 668280
rect 140 667112 633326 667342
rect 0 666771 633326 667112
rect 140 666397 633326 666771
rect 0 666146 633326 666397
rect 140 665916 633326 666146
rect 0 665502 633326 665916
rect 140 665272 633326 665502
rect 0 664858 633326 665272
rect 140 664628 633326 664858
rect 0 664306 633326 664628
rect 140 664076 633326 664306
rect 0 661822 633326 664076
rect 140 661592 633326 661822
rect 0 661178 633326 661592
rect 140 660948 633326 661178
rect 0 660534 633326 660948
rect 140 660304 633326 660534
rect 0 660148 633326 660304
rect 0 659982 633186 660148
rect 140 659926 633186 659982
rect 140 659752 633326 659926
rect 0 658148 633326 659752
rect 0 658142 633186 658148
rect 140 657926 633186 658142
rect 140 657912 633326 657926
rect 0 657498 633326 657912
rect 140 657268 633326 657498
rect 0 656854 633326 657268
rect 140 656624 633186 656854
rect 0 656302 633326 656624
rect 140 656072 633186 656302
rect 0 655658 633326 656072
rect 0 655428 633186 655658
rect 0 655014 633326 655428
rect 0 654784 633186 655014
rect 0 653174 633326 654784
rect 0 652944 633186 653174
rect 0 652622 633326 652944
rect 0 652392 633186 652622
rect 0 651978 633326 652392
rect 0 651748 633186 651978
rect 0 651334 633326 651748
rect 0 651104 633186 651334
rect 0 650784 633326 651104
rect 140 650564 633326 650784
rect 0 648850 633326 650564
rect 0 648784 633186 648850
rect 754 648620 633186 648784
rect 754 648564 633326 648620
rect 0 648298 633326 648564
rect 0 648068 633186 648298
rect 0 647654 633326 648068
rect 0 647424 633186 647654
rect 0 647010 633326 647424
rect 0 646780 633186 647010
rect 0 646529 633326 646780
rect 0 646155 633186 646529
rect 0 645814 633326 646155
rect 0 645584 633186 645814
rect 0 644646 633326 645584
rect 0 644358 633186 644646
rect 0 643974 633326 644358
rect 0 643744 633186 643974
rect 0 642134 633326 643744
rect 0 641904 633186 642134
rect 0 627822 633326 641904
rect 140 627592 633326 627822
rect 0 625982 633326 627592
rect 140 625752 633326 625982
rect 0 625368 633326 625752
rect 140 625080 633326 625368
rect 0 624142 633326 625080
rect 140 623912 633326 624142
rect 0 623571 633326 623912
rect 140 623197 633326 623571
rect 0 622946 633326 623197
rect 140 622716 633326 622946
rect 0 622302 633326 622716
rect 140 622072 633326 622302
rect 0 621658 633326 622072
rect 140 621428 633326 621658
rect 0 621106 633326 621428
rect 140 620876 633326 621106
rect 0 618622 633326 620876
rect 140 618392 633326 618622
rect 0 617978 633326 618392
rect 140 617748 633326 617978
rect 0 617334 633326 617748
rect 140 617104 633326 617334
rect 0 616782 633326 617104
rect 140 616552 633326 616782
rect 0 615148 633326 616552
rect 0 614942 633186 615148
rect 140 614926 633186 614942
rect 140 614712 633326 614926
rect 0 614298 633326 614712
rect 140 614068 633326 614298
rect 0 613654 633326 614068
rect 140 613424 633326 613654
rect 0 613148 633326 613424
rect 0 613102 633186 613148
rect 140 612926 633186 613102
rect 140 612872 633326 612926
rect 0 611654 633326 612872
rect 0 611424 633186 611654
rect 0 611102 633326 611424
rect 0 610872 633186 611102
rect 0 610458 633326 610872
rect 0 610228 633186 610458
rect 0 609814 633326 610228
rect 0 609584 633186 609814
rect 0 607974 633326 609584
rect 0 607784 633186 607974
rect 140 607744 633186 607784
rect 140 607564 633326 607744
rect 0 607422 633326 607564
rect 0 607192 633186 607422
rect 0 606778 633326 607192
rect 0 606548 633186 606778
rect 0 606134 633326 606548
rect 0 605904 633186 606134
rect 0 605784 633326 605904
rect 754 605564 633326 605784
rect 0 603650 633326 605564
rect 0 603420 633186 603650
rect 0 603098 633326 603420
rect 0 602868 633186 603098
rect 0 602454 633326 602868
rect 0 602224 633186 602454
rect 0 601810 633326 602224
rect 0 601580 633186 601810
rect 0 601329 633326 601580
rect 0 600955 633186 601329
rect 0 600614 633326 600955
rect 0 600384 633186 600614
rect 0 599446 633326 600384
rect 0 599158 633186 599446
rect 0 598774 633326 599158
rect 0 598544 633186 598774
rect 0 596934 633326 598544
rect 0 596704 633186 596934
rect 0 584622 633326 596704
rect 140 584392 633326 584622
rect 0 582782 633326 584392
rect 140 582552 633326 582782
rect 0 582168 633326 582552
rect 140 581880 633326 582168
rect 0 580942 633326 581880
rect 140 580712 633326 580942
rect 0 580371 633326 580712
rect 140 579997 633326 580371
rect 0 579746 633326 579997
rect 140 579516 633326 579746
rect 0 579102 633326 579516
rect 140 578872 633326 579102
rect 0 578458 633326 578872
rect 140 578228 633326 578458
rect 0 577906 633326 578228
rect 140 577676 633326 577906
rect 0 575422 633326 577676
rect 140 575192 633326 575422
rect 0 574778 633326 575192
rect 140 574548 633326 574778
rect 0 574134 633326 574548
rect 140 573904 633326 574134
rect 0 573582 633326 573904
rect 140 573352 633326 573582
rect 0 571742 633326 573352
rect 140 571512 633326 571742
rect 0 571098 633326 571512
rect 140 570868 633326 571098
rect 0 570454 633326 570868
rect 140 570224 633326 570454
rect 0 570148 633326 570224
rect 0 569926 633186 570148
rect 0 569902 633326 569926
rect 140 569672 633326 569902
rect 0 568148 633326 569672
rect 0 567926 633186 568148
rect 0 566654 633326 567926
rect 0 566424 633186 566654
rect 0 566102 633326 566424
rect 0 565872 633186 566102
rect 0 565458 633326 565872
rect 0 565228 633186 565458
rect 0 564814 633326 565228
rect 0 564784 633186 564814
rect 140 564584 633186 564784
rect 140 564564 633326 564584
rect 0 562974 633326 564564
rect 0 562784 633186 562974
rect 754 562744 633186 562784
rect 754 562564 633326 562744
rect 0 562422 633326 562564
rect 0 562192 633186 562422
rect 0 561778 633326 562192
rect 0 561548 633186 561778
rect 0 561134 633326 561548
rect 0 560904 633186 561134
rect 0 558650 633326 560904
rect 0 558420 633186 558650
rect 0 558098 633326 558420
rect 0 557868 633186 558098
rect 0 557454 633326 557868
rect 0 557224 633186 557454
rect 0 556810 633326 557224
rect 0 556580 633186 556810
rect 0 556329 633326 556580
rect 0 555955 633186 556329
rect 0 555614 633326 555955
rect 0 555384 633186 555614
rect 0 554446 633326 555384
rect 0 554158 633186 554446
rect 0 553774 633326 554158
rect 0 553544 633186 553774
rect 0 551934 633326 553544
rect 0 551704 633186 551934
rect 0 541422 633326 551704
rect 140 541192 633326 541422
rect 0 539582 633326 541192
rect 140 539352 633326 539582
rect 0 538968 633326 539352
rect 140 538680 633326 538968
rect 0 537742 633326 538680
rect 140 537512 633326 537742
rect 0 537171 633326 537512
rect 140 536797 633326 537171
rect 0 536546 633326 536797
rect 140 536316 633326 536546
rect 0 535902 633326 536316
rect 140 535672 633326 535902
rect 0 535258 633326 535672
rect 140 535028 633326 535258
rect 0 534706 633326 535028
rect 140 534476 633326 534706
rect 0 532222 633326 534476
rect 140 531992 633326 532222
rect 0 531578 633326 531992
rect 140 531348 633326 531578
rect 0 530934 633326 531348
rect 140 530704 633326 530934
rect 0 530382 633326 530704
rect 140 530152 633326 530382
rect 0 528542 633326 530152
rect 140 528312 633326 528542
rect 0 527898 633326 528312
rect 140 527668 633326 527898
rect 0 527254 633326 527668
rect 140 527024 633326 527254
rect 0 526702 633326 527024
rect 140 526472 633326 526702
rect 0 525148 633326 526472
rect 0 524926 633186 525148
rect 0 523147 633326 524926
rect 0 522925 633186 523147
rect 0 521784 633326 522925
rect 140 521564 633326 521784
rect 0 521454 633326 521564
rect 0 521224 633186 521454
rect 0 520902 633326 521224
rect 0 520672 633186 520902
rect 0 520258 633326 520672
rect 0 520028 633186 520258
rect 0 519784 633326 520028
rect 754 519614 633326 519784
rect 754 519564 633186 519614
rect 0 519384 633186 519564
rect 0 517774 633326 519384
rect 0 517544 633186 517774
rect 0 517222 633326 517544
rect 0 516992 633186 517222
rect 0 516578 633326 516992
rect 0 516348 633186 516578
rect 0 515934 633326 516348
rect 0 515704 633186 515934
rect 0 513450 633326 515704
rect 0 513220 633186 513450
rect 0 512898 633326 513220
rect 0 512668 633126 512898
rect 0 512254 633326 512668
rect 0 512024 633186 512254
rect 0 511610 633326 512024
rect 0 511380 633186 511610
rect 0 511129 633326 511380
rect 0 510755 633186 511129
rect 0 510414 633326 510755
rect 0 510184 633186 510414
rect 0 509246 633326 510184
rect 0 508958 633186 509246
rect 0 508574 633326 508958
rect 0 508344 633186 508574
rect 0 506734 633326 508344
rect 0 506504 633186 506734
rect 0 498222 633326 506504
rect 140 497992 633326 498222
rect 0 496382 633326 497992
rect 140 496152 633326 496382
rect 0 495768 633326 496152
rect 140 495480 633326 495768
rect 0 494542 633326 495480
rect 140 494312 633326 494542
rect 0 493971 633326 494312
rect 140 493597 633326 493971
rect 0 493346 633326 493597
rect 140 493116 633326 493346
rect 0 492702 633326 493116
rect 140 492472 633326 492702
rect 0 492058 633326 492472
rect 140 491828 633326 492058
rect 0 491506 633326 491828
rect 140 491276 633326 491506
rect 0 489022 633326 491276
rect 140 488792 633326 489022
rect 0 488378 633326 488792
rect 140 488148 633326 488378
rect 0 487734 633326 488148
rect 140 487504 633326 487734
rect 0 487182 633326 487504
rect 140 486952 633326 487182
rect 0 485342 633326 486952
rect 140 485112 633326 485342
rect 0 484698 633326 485112
rect 140 484468 633326 484698
rect 0 484054 633326 484468
rect 140 483824 633326 484054
rect 0 483502 633326 483824
rect 140 483272 633326 483502
rect 0 478784 633326 483272
rect 140 478564 633326 478784
rect 0 476784 633326 478564
rect 754 476644 633326 476784
rect 754 476564 633186 476644
rect 0 471704 633186 476564
rect 0 466664 633326 471704
rect 0 461724 633186 466664
rect 0 455800 633326 461724
rect 140 450860 633326 455800
rect 0 445822 633326 450860
rect 140 440882 633326 445822
rect 0 432642 633326 440882
rect 0 432562 633186 432642
rect 0 417722 633571 432562
rect 0 417642 633186 417722
rect 0 413684 633326 417642
rect 140 408734 633326 413684
rect 0 408594 633326 408734
rect 140 403782 633326 408594
rect 0 403642 633326 403782
rect 140 398682 633326 403642
rect 0 388444 633326 398682
rect 0 383504 633186 388444
rect 0 378466 633326 383504
rect 0 373526 633186 378466
rect 0 370622 633326 373526
rect 140 370392 633326 370622
rect 0 368782 633326 370392
rect 140 368552 633326 368782
rect 0 368168 633326 368552
rect 140 367880 633326 368168
rect 0 366942 633326 367880
rect 140 366712 633326 366942
rect 0 366371 633326 366712
rect 140 365997 633326 366371
rect 0 365746 633326 365997
rect 140 365516 633326 365746
rect 0 365102 633326 365516
rect 140 364872 633326 365102
rect 0 364458 633326 364872
rect 140 364228 633326 364458
rect 0 363906 633326 364228
rect 140 363676 633326 363906
rect 0 361422 633326 363676
rect 140 361192 633326 361422
rect 0 360778 633326 361192
rect 140 360548 633326 360778
rect 0 360134 633326 360548
rect 140 359904 633326 360134
rect 0 359582 633326 359904
rect 140 359352 633326 359582
rect 0 357742 633326 359352
rect 140 357512 633326 357742
rect 0 357098 633326 357512
rect 140 356868 633326 357098
rect 0 356454 633326 356868
rect 140 356224 633326 356454
rect 0 355902 633326 356224
rect 140 355672 633326 355902
rect 0 349784 633326 355672
rect 140 349564 633326 349784
rect 0 348148 633326 349564
rect 0 347926 633186 348148
rect 0 347784 633326 347926
rect 754 347564 633326 347784
rect 0 346147 633326 347564
rect 0 345925 633186 346147
rect 0 344254 633326 345925
rect 0 344024 633186 344254
rect 0 343702 633326 344024
rect 0 343472 633186 343702
rect 0 343058 633326 343472
rect 0 342828 633186 343058
rect 0 342414 633326 342828
rect 0 342184 633186 342414
rect 0 340574 633326 342184
rect 0 340344 633186 340574
rect 0 340022 633326 340344
rect 0 339792 633186 340022
rect 0 339378 633326 339792
rect 0 339148 633186 339378
rect 0 338734 633326 339148
rect 0 338504 633186 338734
rect 0 336250 633326 338504
rect 0 336020 633186 336250
rect 0 335698 633326 336020
rect 0 335468 633186 335698
rect 0 335054 633326 335468
rect 0 334824 633186 335054
rect 0 334410 633326 334824
rect 0 334180 633186 334410
rect 0 333929 633326 334180
rect 0 333555 633186 333929
rect 0 333214 633326 333555
rect 0 332984 633186 333214
rect 0 332046 633326 332984
rect 0 331758 633186 332046
rect 0 331374 633326 331758
rect 0 331144 633186 331374
rect 0 329534 633326 331144
rect 0 329304 633186 329534
rect 0 327422 633326 329304
rect 140 327192 633326 327422
rect 0 325582 633326 327192
rect 140 325352 633326 325582
rect 0 324968 633326 325352
rect 140 324680 633326 324968
rect 0 323742 633326 324680
rect 140 323512 633326 323742
rect 0 323171 633326 323512
rect 140 322797 633326 323171
rect 0 322546 633326 322797
rect 140 322316 633326 322546
rect 0 321902 633326 322316
rect 140 321672 633326 321902
rect 0 321258 633326 321672
rect 140 321028 633326 321258
rect 0 320706 633326 321028
rect 140 320476 633326 320706
rect 0 318222 633326 320476
rect 140 317992 633326 318222
rect 0 317578 633326 317992
rect 140 317348 633326 317578
rect 0 316934 633326 317348
rect 140 316704 633326 316934
rect 0 316382 633326 316704
rect 140 316152 633326 316382
rect 0 314542 633326 316152
rect 140 314312 633326 314542
rect 0 313898 633326 314312
rect 140 313668 633326 313898
rect 0 313254 633326 313668
rect 140 313024 633326 313254
rect 0 312702 633326 313024
rect 140 312472 633326 312702
rect 0 306784 633326 312472
rect 140 306564 633326 306784
rect 0 304784 633326 306564
rect 754 304564 633326 304784
rect 0 303148 633326 304564
rect 0 302926 633186 303148
rect 0 301147 633326 302926
rect 0 300925 633186 301147
rect 0 299054 633326 300925
rect 0 298824 633186 299054
rect 0 298502 633326 298824
rect 0 298272 633186 298502
rect 0 297858 633326 298272
rect 0 297628 633186 297858
rect 0 297214 633326 297628
rect 0 296984 633186 297214
rect 0 295374 633326 296984
rect 0 295144 633186 295374
rect 0 294822 633326 295144
rect 0 294592 633186 294822
rect 0 294178 633326 294592
rect 0 293948 633186 294178
rect 0 293534 633326 293948
rect 0 293304 633126 293534
rect 0 291050 633326 293304
rect 0 290820 633186 291050
rect 0 290498 633326 290820
rect 0 290268 633186 290498
rect 0 289854 633326 290268
rect 0 289624 633186 289854
rect 0 289210 633326 289624
rect 0 288980 633186 289210
rect 0 288729 633326 288980
rect 0 288355 633186 288729
rect 0 288014 633326 288355
rect 0 287784 633186 288014
rect 0 286846 633326 287784
rect 0 286558 633186 286846
rect 0 286174 633326 286558
rect 0 285944 633186 286174
rect 0 284334 633326 285944
rect 0 284222 633186 284334
rect 140 284104 633186 284222
rect 140 283992 633326 284104
rect 0 282382 633326 283992
rect 140 282152 633326 282382
rect 0 281768 633326 282152
rect 140 281480 633326 281768
rect 0 280542 633326 281480
rect 140 280312 633326 280542
rect 0 279971 633326 280312
rect 140 279597 633326 279971
rect 0 279346 633326 279597
rect 140 279116 633326 279346
rect 0 278702 633326 279116
rect 140 278472 633326 278702
rect 0 278058 633326 278472
rect 140 277828 633326 278058
rect 0 277506 633326 277828
rect 140 277276 633326 277506
rect 0 275022 633326 277276
rect 140 274792 633326 275022
rect 0 274378 633326 274792
rect 140 274148 633326 274378
rect 0 273734 633326 274148
rect 140 273504 633326 273734
rect 0 273182 633326 273504
rect 140 272952 633326 273182
rect 0 271342 633326 272952
rect 140 271112 633326 271342
rect 0 270698 633326 271112
rect 140 270468 633326 270698
rect 0 270054 633326 270468
rect 140 269824 633326 270054
rect 0 269502 633326 269824
rect 140 269272 633326 269502
rect 0 263784 633326 269272
rect 140 263564 633326 263784
rect 0 261784 633326 263564
rect 754 261564 633326 261784
rect 0 258148 633326 261564
rect 0 257926 633186 258148
rect 0 256147 633326 257926
rect 0 255925 633186 256147
rect 0 254054 633326 255925
rect 0 253824 633186 254054
rect 0 253502 633326 253824
rect 0 253272 633186 253502
rect 0 252858 633326 253272
rect 0 252628 633186 252858
rect 0 252214 633326 252628
rect 0 251984 633186 252214
rect 0 250374 633326 251984
rect 0 250144 633186 250374
rect 0 249822 633326 250144
rect 0 249592 633186 249822
rect 0 249178 633326 249592
rect 0 248948 633186 249178
rect 0 248534 633326 248948
rect 0 248304 633186 248534
rect 0 246050 633326 248304
rect 0 245820 633186 246050
rect 0 245498 633326 245820
rect 0 245268 633186 245498
rect 0 244854 633326 245268
rect 0 244624 633186 244854
rect 0 244210 633326 244624
rect 0 243980 633186 244210
rect 0 243729 633326 243980
rect 0 243355 633186 243729
rect 0 243014 633326 243355
rect 0 242784 633186 243014
rect 0 241846 633326 242784
rect 0 241558 633186 241846
rect 0 241174 633326 241558
rect 0 241022 633186 241174
rect 140 240944 633186 241022
rect 140 240792 633326 240944
rect 0 239334 633326 240792
rect 0 239182 633186 239334
rect 140 239104 633186 239182
rect 140 238952 633326 239104
rect 0 238568 633326 238952
rect 140 238280 633326 238568
rect 0 237342 633326 238280
rect 140 237112 633326 237342
rect 0 236771 633326 237112
rect 140 236397 633326 236771
rect 0 236146 633326 236397
rect 140 235916 633326 236146
rect 0 235502 633326 235916
rect 140 235272 633326 235502
rect 0 234858 633326 235272
rect 140 234628 633326 234858
rect 0 234306 633326 234628
rect 140 234076 633326 234306
rect 0 231822 633326 234076
rect 140 231592 633326 231822
rect 0 231178 633326 231592
rect 140 230948 633326 231178
rect 0 230534 633326 230948
rect 140 230304 633326 230534
rect 0 229982 633326 230304
rect 140 229752 633326 229982
rect 0 228142 633326 229752
rect 140 227912 633326 228142
rect 0 227498 633326 227912
rect 140 227268 633326 227498
rect 0 226854 633326 227268
rect 140 226624 633326 226854
rect 0 226302 633326 226624
rect 140 226072 633326 226302
rect 0 220784 633326 226072
rect 140 220564 633326 220784
rect 0 218784 633326 220564
rect 754 218564 633326 218784
rect 0 213148 633326 218564
rect 0 212926 633186 213148
rect 0 211147 633326 212926
rect 0 210925 633186 211147
rect 0 209054 633326 210925
rect 0 208824 633186 209054
rect 0 208502 633326 208824
rect 0 208272 633186 208502
rect 0 207858 633326 208272
rect 0 207628 633186 207858
rect 0 207214 633326 207628
rect 0 206984 633186 207214
rect 0 205374 633326 206984
rect 0 205144 633186 205374
rect 0 204822 633326 205144
rect 0 204592 633186 204822
rect 0 204178 633326 204592
rect 0 203948 633186 204178
rect 0 203534 633326 203948
rect 0 203304 633186 203534
rect 0 201050 633326 203304
rect 0 200820 633186 201050
rect 0 200498 633326 200820
rect 0 200268 633186 200498
rect 0 199854 633326 200268
rect 0 199624 633186 199854
rect 0 199210 633326 199624
rect 0 198980 633186 199210
rect 0 198729 633326 198980
rect 0 198355 633186 198729
rect 0 198014 633326 198355
rect 0 197822 633186 198014
rect 140 197784 633186 197822
rect 140 197592 633326 197784
rect 0 196846 633326 197592
rect 0 196558 633186 196846
rect 0 196174 633326 196558
rect 0 195982 633186 196174
rect 140 195944 633186 195982
rect 140 195752 633326 195944
rect 0 195368 633326 195752
rect 140 195080 633326 195368
rect 0 194334 633326 195080
rect 0 194142 633186 194334
rect 140 194104 633186 194142
rect 140 193912 633326 194104
rect 0 193571 633326 193912
rect 140 193197 633326 193571
rect 0 192946 633326 193197
rect 140 192716 633326 192946
rect 0 192302 633326 192716
rect 140 192072 633326 192302
rect 0 191658 633326 192072
rect 140 191428 633326 191658
rect 0 191106 633326 191428
rect 140 190876 633326 191106
rect 0 188622 633326 190876
rect 140 188392 633326 188622
rect 0 187978 633326 188392
rect 140 187748 633326 187978
rect 0 187334 633326 187748
rect 140 187104 633326 187334
rect 0 186782 633326 187104
rect 140 186552 633326 186782
rect 0 184942 633326 186552
rect 140 184712 633326 184942
rect 0 184298 633326 184712
rect 140 184068 633326 184298
rect 0 183654 633326 184068
rect 140 183424 633326 183654
rect 0 183102 633326 183424
rect 140 182872 633326 183102
rect 0 177784 633326 182872
rect 140 177564 633326 177784
rect 0 175784 633326 177564
rect 754 175564 633326 175784
rect 0 168148 633326 175564
rect 0 167926 633186 168148
rect 0 166147 633326 167926
rect 0 165925 633186 166147
rect 0 163854 633326 165925
rect 0 163624 633186 163854
rect 0 163302 633326 163624
rect 0 163072 633186 163302
rect 0 162658 633326 163072
rect 0 162428 633186 162658
rect 0 162014 633326 162428
rect 0 161784 633186 162014
rect 0 160174 633326 161784
rect 0 159944 633186 160174
rect 0 159622 633326 159944
rect 0 159392 633186 159622
rect 0 158978 633326 159392
rect 0 158748 633186 158978
rect 0 158334 633326 158748
rect 0 158104 633186 158334
rect 0 155850 633326 158104
rect 0 155620 633186 155850
rect 0 155298 633326 155620
rect 0 155068 633186 155298
rect 0 154654 633326 155068
rect 0 154622 633186 154654
rect 140 154424 633186 154622
rect 140 154392 633326 154424
rect 0 154010 633326 154392
rect 0 153780 633186 154010
rect 0 153529 633326 153780
rect 0 153155 633186 153529
rect 0 152814 633326 153155
rect 0 152782 633186 152814
rect 140 152584 633186 152782
rect 140 152552 633326 152584
rect 0 152168 633326 152552
rect 140 151880 633326 152168
rect 0 151646 633326 151880
rect 0 151358 633186 151646
rect 0 150974 633326 151358
rect 0 150942 633186 150974
rect 140 150744 633186 150942
rect 140 150712 633326 150744
rect 0 150371 633326 150712
rect 140 149997 633326 150371
rect 0 149746 633326 149997
rect 140 149516 633326 149746
rect 0 149134 633326 149516
rect 0 149102 633186 149134
rect 140 148904 633186 149102
rect 140 148872 633326 148904
rect 0 148458 633326 148872
rect 140 148228 633326 148458
rect 0 147906 633326 148228
rect 140 147676 633326 147906
rect 0 145422 633326 147676
rect 140 145192 633326 145422
rect 0 144778 633326 145192
rect 140 144548 633326 144778
rect 0 144134 633326 144548
rect 140 143904 633326 144134
rect 0 143582 633326 143904
rect 140 143352 633326 143582
rect 0 141742 633326 143352
rect 140 141512 633326 141742
rect 0 141098 633326 141512
rect 140 140868 633326 141098
rect 0 140454 633326 140868
rect 140 140224 633326 140454
rect 0 139902 633326 140224
rect 140 139672 633326 139902
rect 0 134784 633326 139672
rect 140 134564 633326 134784
rect 0 132784 633326 134564
rect 754 132564 633326 132784
rect 0 123148 633326 132564
rect 0 122926 633186 123148
rect 0 121147 633326 122926
rect 0 120925 633186 121147
rect 0 118854 633326 120925
rect 0 118624 633186 118854
rect 0 118302 633326 118624
rect 0 118072 633186 118302
rect 0 117658 633326 118072
rect 0 117428 633186 117658
rect 0 117014 633326 117428
rect 0 116784 633186 117014
rect 0 115174 633326 116784
rect 0 114944 633186 115174
rect 0 114622 633326 114944
rect 0 114392 633186 114622
rect 0 113978 633326 114392
rect 0 113748 633186 113978
rect 0 113334 633326 113748
rect 0 113104 633186 113334
rect 0 110850 633326 113104
rect 0 110620 633186 110850
rect 0 110298 633326 110620
rect 0 110068 633186 110298
rect 0 109654 633326 110068
rect 0 109424 633186 109654
rect 0 109010 633326 109424
rect 0 108780 633186 109010
rect 0 108529 633326 108780
rect 0 108155 633186 108529
rect 0 107814 633326 108155
rect 0 107584 633186 107814
rect 0 106646 633326 107584
rect 0 106358 633186 106646
rect 0 105974 633326 106358
rect 0 105744 633186 105974
rect 0 104134 633326 105744
rect 0 103904 633186 104134
rect 0 83000 633326 103904
rect 140 78148 633326 83000
rect 140 78060 633186 78148
rect 0 77926 633186 78060
rect 0 76147 633326 77926
rect 0 75925 633186 76147
rect 0 73654 633326 75925
rect 0 73424 633186 73654
rect 0 73102 633326 73424
rect 0 73022 633186 73102
rect 140 72872 633186 73022
rect 140 72458 633326 72872
rect 140 72228 633186 72458
rect 140 71814 633326 72228
rect 140 71584 633186 71814
rect 140 69974 633326 71584
rect 140 69744 633186 69974
rect 140 69422 633326 69744
rect 140 69192 633186 69422
rect 140 68778 633326 69192
rect 140 68548 633186 68778
rect 140 68134 633326 68548
rect 140 68082 633186 68134
rect 0 67904 633186 68082
rect 0 65650 633326 67904
rect 0 65420 633186 65650
rect 0 65098 633326 65420
rect 0 64868 633186 65098
rect 0 64454 633326 64868
rect 0 64224 633186 64454
rect 0 63810 633326 64224
rect 0 63580 633186 63810
rect 0 63329 633326 63580
rect 0 62955 633186 63329
rect 0 62614 633326 62955
rect 0 62384 633186 62614
rect 0 61446 633326 62384
rect 0 61158 633186 61446
rect 0 60774 633326 61158
rect 0 60544 633186 60774
rect 0 58934 633326 60544
rect 0 58704 633186 58934
rect 0 53745 633326 58704
rect 140 53067 633326 53745
rect 0 40884 633326 53067
rect 140 35934 633326 40884
rect 0 30842 633326 35934
rect 140 25882 633326 30842
rect 0 140 633326 25882
rect 0 35 36726 140
rect 41666 35 46704 140
rect 51644 35 199204 140
rect 203994 35 209084 140
rect 214044 35 526926 140
rect 531866 35 536904 140
rect 541844 35 580726 140
rect 585666 35 590704 140
rect 595644 35 633326 140
<< metal4 >>
rect 324 480 4324 952608
rect 4804 4960 8804 948128
rect 11050 480 12330 952608
rect 12970 480 14250 952608
rect 19050 480 20330 952608
rect 20970 480 22250 952608
rect 27050 480 28330 952608
rect 28970 480 30250 952608
rect 35050 480 36330 952608
rect 36970 480 38250 952608
rect 43050 480 44330 952608
rect 44970 480 46250 952608
rect 51050 480 52330 952608
rect 52970 480 54250 952608
rect 59050 480 60330 952608
rect 60970 480 62250 952608
rect 67050 480 68330 952608
rect 68970 480 70250 952608
rect 75050 480 76330 952608
rect 76970 480 78250 952608
rect 83050 480 84330 952608
rect 84970 480 86250 952608
rect 91050 480 92330 952608
rect 92970 480 94250 952608
rect 99050 480 100330 952608
rect 100970 480 102250 952608
rect 107050 480 108330 952608
rect 108970 480 110250 952608
rect 115050 480 116330 952608
rect 116970 480 118250 952608
rect 123050 480 124330 952608
rect 124970 480 126250 952608
rect 131050 480 132330 952608
rect 132970 480 134250 952608
rect 139050 480 140330 952608
rect 140970 480 142250 952608
rect 147050 480 148330 952608
rect 148970 480 150250 952608
rect 155050 480 156330 952608
rect 156970 480 158250 952608
rect 163050 480 164330 952608
rect 164970 480 166250 952608
rect 171050 480 172330 952608
rect 172970 480 174250 952608
rect 179050 480 180330 952608
rect 180970 480 182250 952608
rect 187050 480 188330 952608
rect 188970 480 190250 952608
rect 195050 480 196330 952608
rect 196970 480 198250 952608
rect 203050 480 204330 952608
rect 204970 480 206250 952608
rect 211050 480 212330 952608
rect 212970 480 214250 952608
rect 219050 480 220330 952608
rect 220970 480 222250 952608
rect 227050 480 228330 952608
rect 228970 480 230250 952608
rect 235050 480 236330 952608
rect 236970 480 238250 952608
rect 243050 480 244330 952608
rect 244970 480 246250 952608
rect 251050 480 252330 952608
rect 252970 480 254250 952608
rect 259050 480 260330 952608
rect 260970 480 262250 952608
rect 267050 480 268330 952608
rect 268970 480 270250 952608
rect 275050 480 276330 952608
rect 276970 480 278250 952608
rect 283050 480 284330 952608
rect 284970 480 286250 952608
rect 291050 480 292330 952608
rect 292970 480 294250 952608
rect 299050 480 300330 952608
rect 300970 480 302250 952608
rect 307050 480 308330 952608
rect 308970 480 310250 952608
rect 315050 480 316330 952608
rect 316970 480 318250 952608
rect 323050 480 324330 952608
rect 324970 480 326250 952608
rect 331050 480 332330 952608
rect 332970 480 334250 952608
rect 339050 480 340330 952608
rect 340970 480 342250 952608
rect 347050 480 348330 952608
rect 348970 480 350250 952608
rect 355050 480 356330 952608
rect 356970 480 358250 952608
rect 363050 480 364330 952608
rect 364970 480 366250 952608
rect 371050 480 372330 952608
rect 372970 480 374250 952608
rect 379050 480 380330 952608
rect 380970 480 382250 952608
rect 387050 480 388330 952608
rect 388970 480 390250 952608
rect 395050 480 396330 952608
rect 396970 480 398250 952608
rect 403050 480 404330 952608
rect 404970 480 406250 952608
rect 411050 480 412330 952608
rect 412970 480 414250 952608
rect 419050 480 420330 952608
rect 420970 480 422250 952608
rect 427050 480 428330 952608
rect 428970 480 430250 952608
rect 435050 480 436330 952608
rect 436970 480 438250 952608
rect 443050 480 444330 952608
rect 444970 480 446250 952608
rect 451050 480 452330 952608
rect 452970 480 454250 952608
rect 459050 480 460330 952608
rect 460970 480 462250 952608
rect 467050 480 468330 952608
rect 468970 480 470250 952608
rect 475050 480 476330 952608
rect 476970 480 478250 952608
rect 483050 480 484330 952608
rect 484970 480 486250 952608
rect 491050 480 492330 952608
rect 492970 480 494250 952608
rect 499050 480 500330 952608
rect 500970 480 502250 952608
rect 507050 480 508330 952608
rect 508970 480 510250 952608
rect 515050 480 516330 952608
rect 516970 480 518250 952608
rect 523050 480 524330 952608
rect 524970 480 526250 952608
rect 531050 480 532330 952608
rect 532970 480 534250 952608
rect 539050 480 540330 952608
rect 540970 480 542250 952608
rect 547050 480 548330 952608
rect 548970 480 550250 952608
rect 555050 480 556330 952608
rect 556970 480 558250 952608
rect 563050 480 564330 952608
rect 564970 480 566250 952608
rect 571050 480 572330 952608
rect 572970 480 574250 952608
rect 579050 480 580330 952608
rect 580970 480 582250 952608
rect 587050 480 588330 952608
rect 588970 746596 590250 952608
rect 588970 480 590250 46988
rect 595050 480 596330 952608
rect 596970 480 598250 952608
rect 603050 372861 604330 952608
rect 604970 746596 606250 952608
rect 603050 480 604330 57195
rect 604970 480 606250 46988
rect 611050 480 612330 952608
rect 612970 480 614250 952608
rect 619050 480 620330 952608
rect 620970 480 622250 952608
rect 624524 4960 628524 948128
rect 629004 480 633004 952608
<< obsm4 >>
rect 59 49128 244 922264
rect 4404 49128 4724 922264
rect 8884 49128 10970 922264
rect 12410 49128 12890 922264
rect 14330 49128 18970 922264
rect 20410 49128 20890 922264
rect 22330 49128 26970 922264
rect 28410 49128 28890 922264
rect 30330 49128 34970 922264
rect 36410 49128 36890 922264
rect 38330 49128 42970 922264
rect 44410 49128 44890 922264
rect 46330 49128 50970 922264
rect 52410 49128 52890 922264
rect 54330 49128 58970 922264
rect 60410 49128 60890 922264
rect 62330 49128 66970 922264
rect 68410 49128 68890 922264
rect 70330 49128 74970 922264
rect 76410 49128 76890 922264
rect 78330 49128 82970 922264
rect 84410 49128 84890 922264
rect 86330 49128 90970 922264
rect 92410 49128 92890 922264
rect 94330 49128 98970 922264
rect 100410 49128 100890 922264
rect 102330 49128 106970 922264
rect 108410 49128 108890 922264
rect 110330 49128 114970 922264
rect 116410 49128 116890 922264
rect 118330 49128 122970 922264
rect 124410 49128 124890 922264
rect 126330 49128 130970 922264
rect 132410 49128 132890 922264
rect 134330 49128 138970 922264
rect 140410 49128 140890 922264
rect 142330 49128 146970 922264
rect 148410 49128 148890 922264
rect 150330 49128 154970 922264
rect 156410 49128 156890 922264
rect 158330 49128 162970 922264
rect 164410 49128 164890 922264
rect 166330 49128 170970 922264
rect 172410 49128 172890 922264
rect 174330 49128 178970 922264
rect 180410 49128 180890 922264
rect 182330 49128 186970 922264
rect 188410 49128 188890 922264
rect 190330 49128 194970 922264
rect 196410 49128 196890 922264
rect 198330 49128 202970 922264
rect 204410 49128 204890 922264
rect 206330 49128 210970 922264
rect 212410 49128 212890 922264
rect 214330 49128 218970 922264
rect 220410 49128 220890 922264
rect 222330 49128 226970 922264
rect 228410 49128 228890 922264
rect 230330 49128 234970 922264
rect 236410 49128 236890 922264
rect 238330 49128 242970 922264
rect 244410 49128 244890 922264
rect 246330 49128 250970 922264
rect 252410 49128 252890 922264
rect 254330 49128 258970 922264
rect 260410 49128 260890 922264
rect 262330 49128 266970 922264
rect 268410 49128 268890 922264
rect 270330 49128 274970 922264
rect 276410 49128 276890 922264
rect 278330 49128 282970 922264
rect 284410 49128 284890 922264
rect 286330 49128 290970 922264
rect 292410 49128 292890 922264
rect 294330 49128 298970 922264
rect 300410 49128 300890 922264
rect 302330 49128 306970 922264
rect 308410 49128 308890 922264
rect 310330 49128 314970 922264
rect 316410 49128 316890 922264
rect 318330 49128 322970 922264
rect 324410 49128 324890 922264
rect 326330 49128 330970 922264
rect 332410 49128 332890 922264
rect 334330 49128 338970 922264
rect 340410 49128 340890 922264
rect 342330 49128 346970 922264
rect 348410 49128 348890 922264
rect 350330 49128 354970 922264
rect 356410 49128 356890 922264
rect 358330 49128 362970 922264
rect 364410 49128 364890 922264
rect 366330 49128 370970 922264
rect 372410 49128 372890 922264
rect 374330 49128 378970 922264
rect 380410 49128 380890 922264
rect 382330 49128 386970 922264
rect 388410 49128 388890 922264
rect 390330 49128 394970 922264
rect 396410 49128 396890 922264
rect 398330 49128 402970 922264
rect 404410 49128 404890 922264
rect 406330 49128 410970 922264
rect 412410 49128 412890 922264
rect 414330 49128 418970 922264
rect 420410 49128 420890 922264
rect 422330 49128 426970 922264
rect 428410 49128 428890 922264
rect 430330 49128 434970 922264
rect 436410 49128 436890 922264
rect 438330 49128 442970 922264
rect 444410 49128 444890 922264
rect 446330 49128 450970 922264
rect 452410 49128 452890 922264
rect 454330 49128 458970 922264
rect 460410 49128 460890 922264
rect 462330 49128 466970 922264
rect 468410 49128 468890 922264
rect 470330 49128 474970 922264
rect 476410 49128 476890 922264
rect 478330 49128 482970 922264
rect 484410 49128 484890 922264
rect 486330 49128 490970 922264
rect 492410 49128 492890 922264
rect 494330 49128 498970 922264
rect 500410 49128 500890 922264
rect 502330 49128 506970 922264
rect 508410 49128 508890 922264
rect 510330 49128 514970 922264
rect 516410 49128 516890 922264
rect 518330 49128 522970 922264
rect 524410 49128 524890 922264
rect 526330 49128 530970 922264
rect 532410 49128 532890 922264
rect 534330 49128 538970 922264
rect 540410 49128 540890 922264
rect 542330 49128 546970 922264
rect 548410 49128 548890 922264
rect 550330 49128 554970 922264
rect 556410 49128 556890 922264
rect 558330 49128 562970 922264
rect 564410 49128 564890 922264
rect 566330 49128 570970 922264
rect 572410 49128 572890 922264
rect 574330 49128 578970 922264
rect 580410 49128 580890 922264
rect 582330 49128 586970 922264
rect 588410 746516 588890 922264
rect 590330 746516 594970 922264
rect 588410 49128 594970 746516
rect 596410 49128 596890 922264
rect 598330 372781 602970 922264
rect 604410 746516 604890 922264
rect 606330 746516 610970 922264
rect 604410 372781 610970 746516
rect 598330 57275 610970 372781
rect 598330 49128 602970 57275
rect 604410 49128 610970 57275
rect 612410 49128 612890 922264
rect 614330 49128 618970 922264
rect 620410 49128 620890 922264
rect 622330 49128 624444 922264
rect 628604 49128 628924 922264
rect 633084 49128 633269 922264
<< metal5 >>
rect 324 948608 633004 952608
rect 4804 944128 628524 948128
rect 324 942006 633004 943286
rect 324 940086 633004 941366
rect 324 934006 633004 935286
rect 324 932086 633004 933366
rect 324 926006 633004 927286
rect 324 924086 633004 925366
rect 324 918006 633004 919286
rect 324 916086 633004 917366
rect 324 910006 633004 911286
rect 324 908086 633004 909366
rect 324 902006 633004 903286
rect 324 900086 633004 901366
rect 324 894006 633004 895286
rect 324 892086 633004 893366
rect 324 886006 633004 887286
rect 324 884086 633004 885366
rect 324 878006 633004 879286
rect 324 876086 633004 877366
rect 324 870006 633004 871286
rect 324 868086 633004 869366
rect 324 862006 633004 863286
rect 324 860086 633004 861366
rect 324 854006 633004 855286
rect 324 852086 633004 853366
rect 324 846006 633004 847286
rect 324 844086 633004 845366
rect 324 838006 633004 839286
rect 324 836086 633004 837366
rect 324 830006 633004 831286
rect 324 828086 633004 829366
rect 324 822006 633004 823286
rect 324 820086 633004 821366
rect 324 814006 633004 815286
rect 324 812086 633004 813366
rect 324 806006 633004 807286
rect 324 804086 633004 805366
rect 324 798006 633004 799286
rect 324 796086 633004 797366
rect 324 790006 633004 791286
rect 324 788086 633004 789366
rect 324 782006 633004 783286
rect 324 780086 633004 781366
rect 324 774006 633004 775286
rect 324 772086 633004 773366
rect 324 766006 633004 767286
rect 324 764086 633004 765366
rect 324 758006 633004 759286
rect 324 756086 633004 757366
rect 324 750006 633004 751286
rect 324 748086 633004 749366
rect 324 742006 633004 743286
rect 324 740086 633004 741366
rect 324 734006 633004 735286
rect 324 732086 633004 733366
rect 324 726006 633004 727286
rect 324 724086 633004 725366
rect 324 718006 633004 719286
rect 324 716086 633004 717366
rect 324 710006 633004 711286
rect 324 708086 633004 709366
rect 324 702006 633004 703286
rect 324 700086 633004 701366
rect 324 694006 633004 695286
rect 324 692086 633004 693366
rect 324 686006 633004 687286
rect 324 684086 633004 685366
rect 324 678006 633004 679286
rect 324 676086 633004 677366
rect 324 670006 633004 671286
rect 324 668086 633004 669366
rect 324 662006 633004 663286
rect 324 660086 633004 661366
rect 324 654006 633004 655286
rect 324 652086 633004 653366
rect 324 646006 633004 647286
rect 324 644086 633004 645366
rect 324 638006 633004 639286
rect 324 636086 633004 637366
rect 324 630006 633004 631286
rect 324 628086 633004 629366
rect 324 622006 633004 623286
rect 324 620086 633004 621366
rect 324 614006 633004 615286
rect 324 612086 633004 613366
rect 324 606006 633004 607286
rect 324 604086 633004 605366
rect 324 598006 633004 599286
rect 324 596086 633004 597366
rect 324 590006 633004 591286
rect 324 588086 633004 589366
rect 324 582006 633004 583286
rect 324 580086 633004 581366
rect 324 574006 633004 575286
rect 324 572086 633004 573366
rect 324 566006 633004 567286
rect 324 564086 633004 565366
rect 324 558006 633004 559286
rect 324 556086 633004 557366
rect 324 550006 633004 551286
rect 324 548086 633004 549366
rect 324 542006 633004 543286
rect 324 540086 633004 541366
rect 324 534006 633004 535286
rect 324 532086 633004 533366
rect 324 526006 633004 527286
rect 324 524086 633004 525366
rect 324 518006 633004 519286
rect 324 516086 633004 517366
rect 324 510006 633004 511286
rect 324 508086 633004 509366
rect 324 502006 633004 503286
rect 324 500086 633004 501366
rect 324 494006 633004 495286
rect 324 492086 633004 493366
rect 324 486006 633004 487286
rect 324 484086 633004 485366
rect 324 478006 633004 479286
rect 324 476086 633004 477366
rect 324 470006 633004 471286
rect 324 468086 633004 469366
rect 324 462006 633004 463286
rect 324 460086 633004 461366
rect 324 454006 633004 455286
rect 324 452086 633004 453366
rect 324 446006 633004 447286
rect 324 444086 633004 445366
rect 324 438006 633004 439286
rect 324 436086 633004 437366
rect 324 430006 633004 431286
rect 324 428086 633004 429366
rect 324 422006 633004 423286
rect 324 420086 633004 421366
rect 324 414006 633004 415286
rect 324 412086 633004 413366
rect 324 406006 633004 407286
rect 324 404086 633004 405366
rect 324 398006 633004 399286
rect 324 396086 633004 397366
rect 324 390006 633004 391286
rect 324 388086 633004 389366
rect 324 382006 633004 383286
rect 324 380086 633004 381366
rect 324 374006 633004 375286
rect 324 372086 633004 373366
rect 324 366006 633004 367286
rect 324 364086 633004 365366
rect 324 358006 633004 359286
rect 324 356086 633004 357366
rect 324 350006 633004 351286
rect 324 348086 633004 349366
rect 324 342006 633004 343286
rect 324 340086 633004 341366
rect 324 334006 633004 335286
rect 324 332086 633004 333366
rect 324 326006 633004 327286
rect 324 324086 633004 325366
rect 324 318006 633004 319286
rect 324 316086 633004 317366
rect 324 310006 633004 311286
rect 324 308086 633004 309366
rect 324 302006 633004 303286
rect 324 300086 633004 301366
rect 324 294006 633004 295286
rect 324 292086 633004 293366
rect 324 286006 633004 287286
rect 324 284086 633004 285366
rect 324 278006 633004 279286
rect 324 276086 633004 277366
rect 324 270006 633004 271286
rect 324 268086 633004 269366
rect 324 262006 633004 263286
rect 324 260086 633004 261366
rect 324 254006 633004 255286
rect 324 252086 633004 253366
rect 324 246006 633004 247286
rect 324 244086 633004 245366
rect 324 238006 633004 239286
rect 324 236086 633004 237366
rect 324 230006 633004 231286
rect 324 228086 633004 229366
rect 324 222006 633004 223286
rect 324 220086 633004 221366
rect 324 214006 633004 215286
rect 324 212086 633004 213366
rect 324 206006 633004 207286
rect 324 204086 633004 205366
rect 324 198006 633004 199286
rect 324 196086 633004 197366
rect 324 190006 633004 191286
rect 324 188086 633004 189366
rect 324 182006 633004 183286
rect 324 180086 633004 181366
rect 324 174006 633004 175286
rect 324 172086 633004 173366
rect 324 166006 633004 167286
rect 324 164086 633004 165366
rect 324 158006 633004 159286
rect 324 156086 633004 157366
rect 324 150006 633004 151286
rect 324 148086 633004 149366
rect 324 142006 633004 143286
rect 324 140086 633004 141366
rect 324 134006 633004 135286
rect 324 132086 633004 133366
rect 324 126006 633004 127286
rect 324 124086 633004 125366
rect 324 118006 633004 119286
rect 324 116086 633004 117366
rect 324 110006 633004 111286
rect 324 108086 633004 109366
rect 324 102006 633004 103286
rect 324 100086 633004 101366
rect 324 94006 633004 95286
rect 324 92086 633004 93366
rect 324 86006 633004 87286
rect 324 84086 633004 85366
rect 324 78006 633004 79286
rect 324 76086 633004 77366
rect 324 70006 633004 71286
rect 324 68086 633004 69366
rect 324 62006 633004 63286
rect 324 60086 633004 61366
rect 324 54006 633004 55286
rect 324 52086 633004 53366
rect 324 46006 633004 47286
rect 324 44086 633004 45366
rect 324 38006 633004 39286
rect 324 36086 633004 37366
rect 324 30006 633004 31286
rect 324 28086 633004 29366
rect 324 22006 633004 23286
rect 324 20086 633004 21366
rect 324 14006 633004 15286
rect 324 12086 633004 13366
rect 4804 4960 628524 8960
rect 324 480 633004 4480
<< labels >>
rlabel metal3 s 633266 61238 633726 61366 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 633266 644438 633726 644566 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 633266 689438 633726 689566 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 633266 734438 633726 734566 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 633266 823638 633726 823766 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 633266 912838 633726 912966 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 596360 953270 596488 953726 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 494560 953270 494688 953726 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 443160 953270 443288 953726 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 354160 953270 354288 953726 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 252360 953270 252488 953726 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 633266 106438 633726 106566 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 200760 953270 200888 953726 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 149360 953270 149488 953726 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 97960 953270 98088 953726 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 46560 953270 46688 953726 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -400 924560 60 924688 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -400 754760 60 754888 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -400 711560 60 711688 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -400 668360 60 668488 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -400 625160 60 625288 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s -400 581960 60 582088 4 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 633266 151438 633726 151566 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s -400 538760 60 538888 4 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s -400 495560 60 495688 4 analog_io[31]
port 25 nsew signal bidirectional
rlabel metal3 s -400 367960 60 368088 4 analog_io[32]
port 26 nsew signal bidirectional
rlabel metal3 s -400 324760 60 324888 4 analog_io[33]
port 27 nsew signal bidirectional
rlabel metal3 s -400 281560 60 281688 4 analog_io[34]
port 28 nsew signal bidirectional
rlabel metal3 s -400 238360 60 238488 4 analog_io[35]
port 29 nsew signal bidirectional
rlabel metal3 s -400 195160 60 195288 4 analog_io[36]
port 30 nsew signal bidirectional
rlabel metal3 s -400 151960 60 152088 4 analog_io[37]
port 31 nsew signal bidirectional
rlabel metal2 s 147638 -400 147766 56 8 analog_io[38]
port 32 nsew signal bidirectional
rlabel metal2 s 256238 -400 256366 56 8 analog_io[39]
port 33 nsew signal bidirectional
rlabel metal3 s 633266 196638 633726 196766 6 analog_io[3]
port 34 nsew signal bidirectional
rlabel metal2 s 311038 -400 311166 56 8 analog_io[40]
port 35 nsew signal bidirectional
rlabel metal2 s 365838 -400 365966 56 8 analog_io[41]
port 36 nsew signal bidirectional
rlabel metal2 s 420638 -400 420766 56 8 analog_io[42]
port 37 nsew signal bidirectional
rlabel metal2 s 475438 -400 475566 56 8 analog_io[43]
port 38 nsew signal bidirectional
rlabel metal3 s 633266 241638 633726 241766 6 analog_io[4]
port 39 nsew signal bidirectional
rlabel metal3 s 633266 286638 633726 286766 6 analog_io[5]
port 40 nsew signal bidirectional
rlabel metal3 s 633266 331838 633726 331966 6 analog_io[6]
port 41 nsew signal bidirectional
rlabel metal3 s 633266 509038 633726 509166 6 analog_io[7]
port 42 nsew signal bidirectional
rlabel metal3 s 633266 554238 633726 554366 6 analog_io[8]
port 43 nsew signal bidirectional
rlabel metal3 s 633266 599238 633726 599366 6 analog_io[9]
port 44 nsew signal bidirectional
rlabel metal3 s 633266 63035 633726 63249 6 analog_noesd_io[0]
port 45 nsew signal bidirectional
rlabel metal3 s 633266 646235 633726 646449 6 analog_noesd_io[10]
port 46 nsew signal bidirectional
rlabel metal3 s 633266 691235 633726 691449 6 analog_noesd_io[11]
port 47 nsew signal bidirectional
rlabel metal3 s 633266 736235 633726 736449 6 analog_noesd_io[12]
port 48 nsew signal bidirectional
rlabel metal3 s 633266 825435 633726 825649 6 analog_noesd_io[13]
port 49 nsew signal bidirectional
rlabel metal3 s 633266 914635 633726 914849 6 analog_noesd_io[14]
port 50 nsew signal bidirectional
rlabel metal2 s 594477 953270 594691 953726 6 analog_noesd_io[15]
port 51 nsew signal bidirectional
rlabel metal2 s 492677 953270 492891 953726 6 analog_noesd_io[16]
port 52 nsew signal bidirectional
rlabel metal2 s 441277 953270 441491 953726 6 analog_noesd_io[17]
port 53 nsew signal bidirectional
rlabel metal2 s 352277 953270 352491 953726 6 analog_noesd_io[18]
port 54 nsew signal bidirectional
rlabel metal2 s 250477 953270 250691 953726 6 analog_noesd_io[19]
port 55 nsew signal bidirectional
rlabel metal3 s 633266 108235 633726 108449 6 analog_noesd_io[1]
port 56 nsew signal bidirectional
rlabel metal2 s 198877 953270 199091 953726 6 analog_noesd_io[20]
port 57 nsew signal bidirectional
rlabel metal2 s 147477 953270 147691 953726 6 analog_noesd_io[21]
port 58 nsew signal bidirectional
rlabel metal2 s 96077 953270 96291 953726 6 analog_noesd_io[22]
port 59 nsew signal bidirectional
rlabel metal2 s 44677 953270 44891 953726 6 analog_noesd_io[23]
port 60 nsew signal bidirectional
rlabel metal3 s -400 922677 60 922891 4 analog_noesd_io[24]
port 61 nsew signal bidirectional
rlabel metal3 s -400 752877 60 753091 4 analog_noesd_io[25]
port 62 nsew signal bidirectional
rlabel metal3 s -400 709677 60 709891 4 analog_noesd_io[26]
port 63 nsew signal bidirectional
rlabel metal3 s -400 666477 60 666691 4 analog_noesd_io[27]
port 64 nsew signal bidirectional
rlabel metal3 s -400 623277 60 623491 4 analog_noesd_io[28]
port 65 nsew signal bidirectional
rlabel metal3 s -400 580077 60 580291 4 analog_noesd_io[29]
port 66 nsew signal bidirectional
rlabel metal3 s 633266 153235 633726 153449 6 analog_noesd_io[2]
port 67 nsew signal bidirectional
rlabel metal3 s -400 536877 60 537091 4 analog_noesd_io[30]
port 68 nsew signal bidirectional
rlabel metal3 s -400 493677 60 493891 4 analog_noesd_io[31]
port 69 nsew signal bidirectional
rlabel metal3 s -400 366077 60 366291 4 analog_noesd_io[32]
port 70 nsew signal bidirectional
rlabel metal3 s -400 322877 60 323091 4 analog_noesd_io[33]
port 71 nsew signal bidirectional
rlabel metal3 s -400 279677 60 279891 4 analog_noesd_io[34]
port 72 nsew signal bidirectional
rlabel metal3 s -400 236477 60 236691 4 analog_noesd_io[35]
port 73 nsew signal bidirectional
rlabel metal3 s -400 193277 60 193491 4 analog_noesd_io[36]
port 74 nsew signal bidirectional
rlabel metal3 s -400 150077 60 150291 4 analog_noesd_io[37]
port 75 nsew signal bidirectional
rlabel metal2 s 149435 -400 149649 56 8 analog_noesd_io[38]
port 76 nsew signal bidirectional
rlabel metal2 s 258035 -400 258249 56 8 analog_noesd_io[39]
port 77 nsew signal bidirectional
rlabel metal3 s 633266 198435 633726 198649 6 analog_noesd_io[3]
port 78 nsew signal bidirectional
rlabel metal2 s 312835 -400 313049 56 8 analog_noesd_io[40]
port 79 nsew signal bidirectional
rlabel metal2 s 367635 -400 367849 56 8 analog_noesd_io[41]
port 80 nsew signal bidirectional
rlabel metal2 s 422435 -400 422649 56 8 analog_noesd_io[42]
port 81 nsew signal bidirectional
rlabel metal2 s 477235 -400 477449 56 8 analog_noesd_io[43]
port 82 nsew signal bidirectional
rlabel metal3 s 633266 243435 633726 243649 6 analog_noesd_io[4]
port 83 nsew signal bidirectional
rlabel metal3 s 633266 288435 633726 288649 6 analog_noesd_io[5]
port 84 nsew signal bidirectional
rlabel metal3 s 633266 333635 633726 333849 6 analog_noesd_io[6]
port 85 nsew signal bidirectional
rlabel metal3 s 633266 510835 633726 511049 6 analog_noesd_io[7]
port 86 nsew signal bidirectional
rlabel metal3 s 633266 556035 633726 556249 6 analog_noesd_io[8]
port 87 nsew signal bidirectional
rlabel metal3 s 633266 601035 633726 601249 6 analog_noesd_io[9]
port 88 nsew signal bidirectional
rlabel metal3 s 633266 63660 633726 63730 6 gpio_analog_en[0]
port 89 nsew signal output
rlabel metal3 s 633266 646860 633726 646930 6 gpio_analog_en[10]
port 90 nsew signal output
rlabel metal3 s 633266 691860 633726 691930 6 gpio_analog_en[11]
port 91 nsew signal output
rlabel metal3 s 633266 736860 633726 736930 6 gpio_analog_en[12]
port 92 nsew signal output
rlabel metal3 s 633266 826060 633726 826130 6 gpio_analog_en[13]
port 93 nsew signal output
rlabel metal3 s 633266 915260 633726 915330 6 gpio_analog_en[14]
port 94 nsew signal output
rlabel metal2 s 594004 953270 594060 953726 6 gpio_analog_en[15]
port 95 nsew signal output
rlabel metal2 s 492204 953270 492260 953726 6 gpio_analog_en[16]
port 96 nsew signal output
rlabel metal2 s 440804 953270 440860 953726 6 gpio_analog_en[17]
port 97 nsew signal output
rlabel metal2 s 351804 953270 351860 953726 6 gpio_analog_en[18]
port 98 nsew signal output
rlabel metal2 s 250004 953270 250060 953726 6 gpio_analog_en[19]
port 99 nsew signal output
rlabel metal3 s 633266 108860 633726 108930 6 gpio_analog_en[1]
port 100 nsew signal output
rlabel metal2 s 198404 953270 198460 953726 6 gpio_analog_en[20]
port 101 nsew signal output
rlabel metal2 s 147004 953270 147060 953726 6 gpio_analog_en[21]
port 102 nsew signal output
rlabel metal2 s 95604 953270 95660 953726 6 gpio_analog_en[22]
port 103 nsew signal output
rlabel metal2 s 44204 953270 44260 953726 6 gpio_analog_en[23]
port 104 nsew signal output
rlabel metal3 s -400 922196 60 922266 4 gpio_analog_en[24]
port 105 nsew signal output
rlabel metal3 s -400 752396 60 752466 4 gpio_analog_en[25]
port 106 nsew signal output
rlabel metal3 s -400 709196 60 709266 4 gpio_analog_en[26]
port 107 nsew signal output
rlabel metal3 s -400 665996 60 666066 4 gpio_analog_en[27]
port 108 nsew signal output
rlabel metal3 s -400 622796 60 622866 4 gpio_analog_en[28]
port 109 nsew signal output
rlabel metal3 s -400 579596 60 579666 4 gpio_analog_en[29]
port 110 nsew signal output
rlabel metal3 s 633266 153860 633726 153930 6 gpio_analog_en[2]
port 111 nsew signal output
rlabel metal3 s -400 536396 60 536466 4 gpio_analog_en[30]
port 112 nsew signal output
rlabel metal3 s -400 493196 60 493266 4 gpio_analog_en[31]
port 113 nsew signal output
rlabel metal3 s -400 365596 60 365666 4 gpio_analog_en[32]
port 114 nsew signal output
rlabel metal3 s -400 322396 60 322466 4 gpio_analog_en[33]
port 115 nsew signal output
rlabel metal3 s -400 279196 60 279266 4 gpio_analog_en[34]
port 116 nsew signal output
rlabel metal3 s -400 235996 60 236066 4 gpio_analog_en[35]
port 117 nsew signal output
rlabel metal3 s -400 192796 60 192866 4 gpio_analog_en[36]
port 118 nsew signal output
rlabel metal3 s -400 149596 60 149666 4 gpio_analog_en[37]
port 119 nsew signal output
rlabel metal2 s 150066 -400 150122 56 8 gpio_analog_en[38]
port 120 nsew signal output
rlabel metal2 s 258666 -400 258722 56 8 gpio_analog_en[39]
port 121 nsew signal output
rlabel metal3 s 633266 199060 633726 199130 6 gpio_analog_en[3]
port 122 nsew signal output
rlabel metal2 s 313466 -400 313522 56 8 gpio_analog_en[40]
port 123 nsew signal output
rlabel metal2 s 368266 -400 368322 56 8 gpio_analog_en[41]
port 124 nsew signal output
rlabel metal2 s 423066 -400 423122 56 8 gpio_analog_en[42]
port 125 nsew signal output
rlabel metal2 s 477866 -400 477922 56 8 gpio_analog_en[43]
port 126 nsew signal output
rlabel metal3 s 633266 244060 633726 244130 6 gpio_analog_en[4]
port 127 nsew signal output
rlabel metal3 s 633266 289060 633726 289130 6 gpio_analog_en[5]
port 128 nsew signal output
rlabel metal3 s 633266 334260 633726 334330 6 gpio_analog_en[6]
port 129 nsew signal output
rlabel metal3 s 633266 511460 633726 511530 6 gpio_analog_en[7]
port 130 nsew signal output
rlabel metal3 s 633266 556660 633726 556730 6 gpio_analog_en[8]
port 131 nsew signal output
rlabel metal3 s 633266 601660 633726 601730 6 gpio_analog_en[9]
port 132 nsew signal output
rlabel metal3 s 633266 64948 633726 65018 6 gpio_analog_pol[0]
port 133 nsew signal output
rlabel metal3 s 633266 648148 633726 648218 6 gpio_analog_pol[10]
port 134 nsew signal output
rlabel metal3 s 633266 693148 633726 693218 6 gpio_analog_pol[11]
port 135 nsew signal output
rlabel metal3 s 633266 738148 633726 738218 6 gpio_analog_pol[12]
port 136 nsew signal output
rlabel metal3 s 633266 827348 633726 827418 6 gpio_analog_pol[13]
port 137 nsew signal output
rlabel metal3 s 633266 916548 633726 916618 6 gpio_analog_pol[14]
port 138 nsew signal output
rlabel metal2 s 592716 953270 592772 953726 6 gpio_analog_pol[15]
port 139 nsew signal output
rlabel metal2 s 490916 953270 490972 953726 6 gpio_analog_pol[16]
port 140 nsew signal output
rlabel metal2 s 439516 953270 439572 953726 6 gpio_analog_pol[17]
port 141 nsew signal output
rlabel metal2 s 350516 953270 350572 953726 6 gpio_analog_pol[18]
port 142 nsew signal output
rlabel metal2 s 248716 953270 248772 953726 6 gpio_analog_pol[19]
port 143 nsew signal output
rlabel metal3 s 633266 110148 633726 110218 6 gpio_analog_pol[1]
port 144 nsew signal output
rlabel metal2 s 197116 953270 197172 953726 6 gpio_analog_pol[20]
port 145 nsew signal output
rlabel metal2 s 145716 953244 145772 953726 6 gpio_analog_pol[21]
port 146 nsew signal output
rlabel metal2 s 94316 953270 94372 953726 6 gpio_analog_pol[22]
port 147 nsew signal output
rlabel metal2 s 42916 953270 42972 953726 6 gpio_analog_pol[23]
port 148 nsew signal output
rlabel metal3 s -400 920908 60 920978 4 gpio_analog_pol[24]
port 149 nsew signal output
rlabel metal3 s -400 751108 60 751178 4 gpio_analog_pol[25]
port 150 nsew signal output
rlabel metal3 s -400 707908 60 707978 4 gpio_analog_pol[26]
port 151 nsew signal output
rlabel metal3 s -400 664708 60 664778 4 gpio_analog_pol[27]
port 152 nsew signal output
rlabel metal3 s -400 621508 60 621578 4 gpio_analog_pol[28]
port 153 nsew signal output
rlabel metal3 s -400 578308 60 578378 4 gpio_analog_pol[29]
port 154 nsew signal output
rlabel metal3 s 633266 155148 633726 155218 6 gpio_analog_pol[2]
port 155 nsew signal output
rlabel metal3 s -400 535108 60 535178 4 gpio_analog_pol[30]
port 156 nsew signal output
rlabel metal3 s -400 491908 60 491978 4 gpio_analog_pol[31]
port 157 nsew signal output
rlabel metal3 s -400 364308 60 364378 4 gpio_analog_pol[32]
port 158 nsew signal output
rlabel metal3 s -400 321108 60 321178 4 gpio_analog_pol[33]
port 159 nsew signal output
rlabel metal3 s -400 277908 60 277978 4 gpio_analog_pol[34]
port 160 nsew signal output
rlabel metal3 s -400 234708 60 234778 4 gpio_analog_pol[35]
port 161 nsew signal output
rlabel metal3 s -400 191508 60 191578 4 gpio_analog_pol[36]
port 162 nsew signal output
rlabel metal3 s -400 148308 60 148378 4 gpio_analog_pol[37]
port 163 nsew signal output
rlabel metal2 s 151354 -400 151410 56 8 gpio_analog_pol[38]
port 164 nsew signal output
rlabel metal2 s 259954 -400 260010 56 8 gpio_analog_pol[39]
port 165 nsew signal output
rlabel metal3 s 633266 200348 633726 200418 6 gpio_analog_pol[3]
port 166 nsew signal output
rlabel metal2 s 314754 -400 314810 56 8 gpio_analog_pol[40]
port 167 nsew signal output
rlabel metal2 s 369554 -400 369610 56 8 gpio_analog_pol[41]
port 168 nsew signal output
rlabel metal2 s 424354 -400 424410 56 8 gpio_analog_pol[42]
port 169 nsew signal output
rlabel metal2 s 479154 -400 479210 56 8 gpio_analog_pol[43]
port 170 nsew signal output
rlabel metal3 s 633266 245348 633726 245418 6 gpio_analog_pol[4]
port 171 nsew signal output
rlabel metal3 s 633266 290348 633726 290418 6 gpio_analog_pol[5]
port 172 nsew signal output
rlabel metal3 s 633266 335548 633726 335618 6 gpio_analog_pol[6]
port 173 nsew signal output
rlabel metal3 s 633206 512748 633726 512818 6 gpio_analog_pol[7]
port 174 nsew signal output
rlabel metal3 s 633266 557948 633726 558018 6 gpio_analog_pol[8]
port 175 nsew signal output
rlabel metal3 s 633266 602948 633726 603018 6 gpio_analog_pol[9]
port 176 nsew signal output
rlabel metal3 s 633266 67984 633726 68054 6 gpio_analog_sel[0]
port 177 nsew signal output
rlabel metal3 s 633266 651184 633726 651254 6 gpio_analog_sel[10]
port 178 nsew signal output
rlabel metal3 s 633266 696184 633726 696254 6 gpio_analog_sel[11]
port 179 nsew signal output
rlabel metal3 s 633206 741184 633726 741254 6 gpio_analog_sel[12]
port 180 nsew signal output
rlabel metal3 s 633266 830384 633726 830454 6 gpio_analog_sel[13]
port 181 nsew signal output
rlabel metal3 s 633266 919584 633726 919654 6 gpio_analog_sel[14]
port 182 nsew signal output
rlabel metal2 s 589680 953270 589736 953726 6 gpio_analog_sel[15]
port 183 nsew signal output
rlabel metal2 s 487880 953270 487936 953726 6 gpio_analog_sel[16]
port 184 nsew signal output
rlabel metal2 s 436480 953270 436536 953726 6 gpio_analog_sel[17]
port 185 nsew signal output
rlabel metal2 s 347480 953270 347536 953726 6 gpio_analog_sel[18]
port 186 nsew signal output
rlabel metal2 s 245680 953244 245736 953726 6 gpio_analog_sel[19]
port 187 nsew signal output
rlabel metal3 s 633266 113184 633726 113254 6 gpio_analog_sel[1]
port 188 nsew signal output
rlabel metal2 s 194080 953270 194136 953726 6 gpio_analog_sel[20]
port 189 nsew signal output
rlabel metal2 s 142680 953270 142736 953726 6 gpio_analog_sel[21]
port 190 nsew signal output
rlabel metal2 s 91280 953270 91336 953726 6 gpio_analog_sel[22]
port 191 nsew signal output
rlabel metal2 s 39880 953270 39936 953726 6 gpio_analog_sel[23]
port 192 nsew signal output
rlabel metal3 s -400 917872 60 917942 4 gpio_analog_sel[24]
port 193 nsew signal output
rlabel metal3 s -400 748072 60 748142 4 gpio_analog_sel[25]
port 194 nsew signal output
rlabel metal3 s -400 704872 60 704942 4 gpio_analog_sel[26]
port 195 nsew signal output
rlabel metal3 s -400 661672 60 661742 4 gpio_analog_sel[27]
port 196 nsew signal output
rlabel metal3 s -400 618472 60 618542 4 gpio_analog_sel[28]
port 197 nsew signal output
rlabel metal3 s -400 575272 60 575342 4 gpio_analog_sel[29]
port 198 nsew signal output
rlabel metal3 s 633266 158184 633726 158254 6 gpio_analog_sel[2]
port 199 nsew signal output
rlabel metal3 s -400 532072 60 532142 4 gpio_analog_sel[30]
port 200 nsew signal output
rlabel metal3 s -400 488872 60 488942 4 gpio_analog_sel[31]
port 201 nsew signal output
rlabel metal3 s -400 361272 60 361342 4 gpio_analog_sel[32]
port 202 nsew signal output
rlabel metal3 s -400 318072 60 318142 4 gpio_analog_sel[33]
port 203 nsew signal output
rlabel metal3 s -400 274872 60 274942 4 gpio_analog_sel[34]
port 204 nsew signal output
rlabel metal3 s -400 231672 60 231742 4 gpio_analog_sel[35]
port 205 nsew signal output
rlabel metal3 s -400 188472 60 188542 4 gpio_analog_sel[36]
port 206 nsew signal output
rlabel metal3 s -400 145272 60 145342 4 gpio_analog_sel[37]
port 207 nsew signal output
rlabel metal2 s 154390 -400 154446 56 8 gpio_analog_sel[38]
port 208 nsew signal output
rlabel metal2 s 262990 -400 263046 56 8 gpio_analog_sel[39]
port 209 nsew signal output
rlabel metal3 s 633266 203384 633726 203454 6 gpio_analog_sel[3]
port 210 nsew signal output
rlabel metal2 s 317790 -400 317846 56 8 gpio_analog_sel[40]
port 211 nsew signal output
rlabel metal2 s 372590 -400 372646 56 8 gpio_analog_sel[41]
port 212 nsew signal output
rlabel metal2 s 427390 -400 427446 56 8 gpio_analog_sel[42]
port 213 nsew signal output
rlabel metal2 s 482190 -400 482246 56 8 gpio_analog_sel[43]
port 214 nsew signal output
rlabel metal3 s 633266 248384 633726 248454 6 gpio_analog_sel[4]
port 215 nsew signal output
rlabel metal3 s 633206 293384 633726 293454 6 gpio_analog_sel[5]
port 216 nsew signal output
rlabel metal3 s 633266 338584 633726 338654 6 gpio_analog_sel[6]
port 217 nsew signal output
rlabel metal3 s 633266 515784 633726 515854 6 gpio_analog_sel[7]
port 218 nsew signal output
rlabel metal3 s 633266 560984 633726 561054 6 gpio_analog_sel[8]
port 219 nsew signal output
rlabel metal3 s 633266 605984 633726 606054 6 gpio_analog_sel[9]
port 220 nsew signal output
rlabel metal3 s 633266 64304 633726 64374 6 gpio_dm0[0]
port 221 nsew signal output
rlabel metal3 s 633266 647504 633726 647574 6 gpio_dm0[10]
port 222 nsew signal output
rlabel metal3 s 633266 692504 633726 692574 6 gpio_dm0[11]
port 223 nsew signal output
rlabel metal3 s 633266 737504 633726 737574 6 gpio_dm0[12]
port 224 nsew signal output
rlabel metal3 s 633266 826704 633726 826774 6 gpio_dm0[13]
port 225 nsew signal output
rlabel metal3 s 633266 915904 633726 915974 6 gpio_dm0[14]
port 226 nsew signal output
rlabel metal2 s 593360 953270 593416 953726 6 gpio_dm0[15]
port 227 nsew signal output
rlabel metal2 s 491560 953270 491616 953726 6 gpio_dm0[16]
port 228 nsew signal output
rlabel metal2 s 440160 953270 440216 953726 6 gpio_dm0[17]
port 229 nsew signal output
rlabel metal2 s 351160 953270 351216 953726 6 gpio_dm0[18]
port 230 nsew signal output
rlabel metal2 s 249360 953270 249416 953726 6 gpio_dm0[19]
port 231 nsew signal output
rlabel metal3 s 633266 109504 633726 109574 6 gpio_dm0[1]
port 232 nsew signal output
rlabel metal2 s 197760 953270 197816 953726 6 gpio_dm0[20]
port 233 nsew signal output
rlabel metal2 s 146360 953270 146416 953726 6 gpio_dm0[21]
port 234 nsew signal output
rlabel metal2 s 94960 953270 95016 953726 6 gpio_dm0[22]
port 235 nsew signal output
rlabel metal2 s 43560 953270 43616 953726 6 gpio_dm0[23]
port 236 nsew signal output
rlabel metal3 s -400 921552 60 921622 4 gpio_dm0[24]
port 237 nsew signal output
rlabel metal3 s -400 751752 60 751822 4 gpio_dm0[25]
port 238 nsew signal output
rlabel metal3 s -400 708552 60 708622 4 gpio_dm0[26]
port 239 nsew signal output
rlabel metal3 s -400 665352 60 665422 4 gpio_dm0[27]
port 240 nsew signal output
rlabel metal3 s -400 622152 60 622222 4 gpio_dm0[28]
port 241 nsew signal output
rlabel metal3 s -400 578952 60 579022 4 gpio_dm0[29]
port 242 nsew signal output
rlabel metal3 s 633266 154504 633726 154574 6 gpio_dm0[2]
port 243 nsew signal output
rlabel metal3 s -400 535752 60 535822 4 gpio_dm0[30]
port 244 nsew signal output
rlabel metal3 s -400 492552 60 492622 4 gpio_dm0[31]
port 245 nsew signal output
rlabel metal3 s -400 364952 60 365022 4 gpio_dm0[32]
port 246 nsew signal output
rlabel metal3 s -400 321752 60 321822 4 gpio_dm0[33]
port 247 nsew signal output
rlabel metal3 s -400 278552 60 278622 4 gpio_dm0[34]
port 248 nsew signal output
rlabel metal3 s -400 235352 60 235422 4 gpio_dm0[35]
port 249 nsew signal output
rlabel metal3 s -400 192152 60 192222 4 gpio_dm0[36]
port 250 nsew signal output
rlabel metal3 s -400 148952 60 149022 4 gpio_dm0[37]
port 251 nsew signal output
rlabel metal2 s 150710 -400 150766 56 8 gpio_dm0[38]
port 252 nsew signal output
rlabel metal2 s 259310 -400 259366 56 8 gpio_dm0[39]
port 253 nsew signal output
rlabel metal3 s 633266 199704 633726 199774 6 gpio_dm0[3]
port 254 nsew signal output
rlabel metal2 s 314110 -400 314166 56 8 gpio_dm0[40]
port 255 nsew signal output
rlabel metal2 s 368910 -400 368966 56 8 gpio_dm0[41]
port 256 nsew signal output
rlabel metal2 s 423710 -400 423766 56 8 gpio_dm0[42]
port 257 nsew signal output
rlabel metal2 s 478510 -400 478566 56 8 gpio_dm0[43]
port 258 nsew signal output
rlabel metal3 s 633266 244704 633726 244774 6 gpio_dm0[4]
port 259 nsew signal output
rlabel metal3 s 633266 289704 633726 289774 6 gpio_dm0[5]
port 260 nsew signal output
rlabel metal3 s 633266 334904 633726 334974 6 gpio_dm0[6]
port 261 nsew signal output
rlabel metal3 s 633266 512104 633726 512174 6 gpio_dm0[7]
port 262 nsew signal output
rlabel metal3 s 633266 557304 633726 557374 6 gpio_dm0[8]
port 263 nsew signal output
rlabel metal3 s 633266 602304 633726 602374 6 gpio_dm0[9]
port 264 nsew signal output
rlabel metal3 s 633266 62464 633726 62534 6 gpio_dm1[0]
port 265 nsew signal output
rlabel metal3 s 633266 645664 633726 645734 6 gpio_dm1[10]
port 266 nsew signal output
rlabel metal3 s 633266 690664 633726 690734 6 gpio_dm1[11]
port 267 nsew signal output
rlabel metal3 s 633266 735664 633726 735734 6 gpio_dm1[12]
port 268 nsew signal output
rlabel metal3 s 633266 824864 633726 824934 6 gpio_dm1[13]
port 269 nsew signal output
rlabel metal3 s 633266 914064 633726 914134 6 gpio_dm1[14]
port 270 nsew signal output
rlabel metal2 s 595200 953270 595256 953726 6 gpio_dm1[15]
port 271 nsew signal output
rlabel metal2 s 493400 953270 493456 953726 6 gpio_dm1[16]
port 272 nsew signal output
rlabel metal2 s 442000 953270 442056 953726 6 gpio_dm1[17]
port 273 nsew signal output
rlabel metal2 s 353000 953270 353056 953726 6 gpio_dm1[18]
port 274 nsew signal output
rlabel metal2 s 251200 953270 251256 953726 6 gpio_dm1[19]
port 275 nsew signal output
rlabel metal3 s 633266 107664 633726 107734 6 gpio_dm1[1]
port 276 nsew signal output
rlabel metal2 s 199600 953270 199656 953726 6 gpio_dm1[20]
port 277 nsew signal output
rlabel metal2 s 148200 953270 148256 953726 6 gpio_dm1[21]
port 278 nsew signal output
rlabel metal2 s 96800 953270 96856 953726 6 gpio_dm1[22]
port 279 nsew signal output
rlabel metal2 s 45400 953270 45456 953726 6 gpio_dm1[23]
port 280 nsew signal output
rlabel metal3 s -400 923392 60 923462 4 gpio_dm1[24]
port 281 nsew signal output
rlabel metal3 s -400 753592 60 753662 4 gpio_dm1[25]
port 282 nsew signal output
rlabel metal3 s -400 710392 60 710462 4 gpio_dm1[26]
port 283 nsew signal output
rlabel metal3 s -400 667192 60 667262 4 gpio_dm1[27]
port 284 nsew signal output
rlabel metal3 s -400 623992 60 624062 4 gpio_dm1[28]
port 285 nsew signal output
rlabel metal3 s -400 580792 60 580862 4 gpio_dm1[29]
port 286 nsew signal output
rlabel metal3 s 633266 152664 633726 152734 6 gpio_dm1[2]
port 287 nsew signal output
rlabel metal3 s -400 537592 60 537662 4 gpio_dm1[30]
port 288 nsew signal output
rlabel metal3 s -400 494392 60 494462 4 gpio_dm1[31]
port 289 nsew signal output
rlabel metal3 s -400 366792 60 366862 4 gpio_dm1[32]
port 290 nsew signal output
rlabel metal3 s -400 323592 60 323662 4 gpio_dm1[33]
port 291 nsew signal output
rlabel metal3 s -400 280392 60 280462 4 gpio_dm1[34]
port 292 nsew signal output
rlabel metal3 s -400 237192 60 237262 4 gpio_dm1[35]
port 293 nsew signal output
rlabel metal3 s -400 193992 60 194062 4 gpio_dm1[36]
port 294 nsew signal output
rlabel metal3 s -400 150792 60 150862 4 gpio_dm1[37]
port 295 nsew signal output
rlabel metal2 s 148870 -400 148926 56 8 gpio_dm1[38]
port 296 nsew signal output
rlabel metal2 s 257470 -400 257526 56 8 gpio_dm1[39]
port 297 nsew signal output
rlabel metal3 s 633266 197864 633726 197934 6 gpio_dm1[3]
port 298 nsew signal output
rlabel metal2 s 312270 -400 312326 56 8 gpio_dm1[40]
port 299 nsew signal output
rlabel metal2 s 367070 -400 367126 56 8 gpio_dm1[41]
port 300 nsew signal output
rlabel metal2 s 421870 -400 421926 56 8 gpio_dm1[42]
port 301 nsew signal output
rlabel metal2 s 476670 -400 476726 56 8 gpio_dm1[43]
port 302 nsew signal output
rlabel metal3 s 633266 242864 633726 242934 6 gpio_dm1[4]
port 303 nsew signal output
rlabel metal3 s 633266 287864 633726 287934 6 gpio_dm1[5]
port 304 nsew signal output
rlabel metal3 s 633266 333064 633726 333134 6 gpio_dm1[6]
port 305 nsew signal output
rlabel metal3 s 633266 510264 633726 510334 6 gpio_dm1[7]
port 306 nsew signal output
rlabel metal3 s 633266 555464 633726 555534 6 gpio_dm1[8]
port 307 nsew signal output
rlabel metal3 s 633266 600464 633726 600534 6 gpio_dm1[9]
port 308 nsew signal output
rlabel metal3 s 633266 68628 633726 68698 6 gpio_dm2[0]
port 309 nsew signal output
rlabel metal3 s 633266 651828 633726 651898 6 gpio_dm2[10]
port 310 nsew signal output
rlabel metal3 s 633266 696828 633726 696898 6 gpio_dm2[11]
port 311 nsew signal output
rlabel metal3 s 633266 741828 633726 741898 6 gpio_dm2[12]
port 312 nsew signal output
rlabel metal3 s 633266 831028 633726 831098 6 gpio_dm2[13]
port 313 nsew signal output
rlabel metal3 s 633266 920228 633726 920298 6 gpio_dm2[14]
port 314 nsew signal output
rlabel metal2 s 589036 953270 589092 953726 6 gpio_dm2[15]
port 315 nsew signal output
rlabel metal2 s 487236 953270 487292 953726 6 gpio_dm2[16]
port 316 nsew signal output
rlabel metal2 s 435836 953270 435892 953726 6 gpio_dm2[17]
port 317 nsew signal output
rlabel metal2 s 346836 953270 346892 953726 6 gpio_dm2[18]
port 318 nsew signal output
rlabel metal2 s 245036 953270 245092 953726 6 gpio_dm2[19]
port 319 nsew signal output
rlabel metal3 s 633266 113828 633726 113898 6 gpio_dm2[1]
port 320 nsew signal output
rlabel metal2 s 193436 953270 193492 953726 6 gpio_dm2[20]
port 321 nsew signal output
rlabel metal2 s 142036 953270 142092 953726 6 gpio_dm2[21]
port 322 nsew signal output
rlabel metal2 s 90636 953270 90692 953726 6 gpio_dm2[22]
port 323 nsew signal output
rlabel metal2 s 39236 953270 39292 953726 6 gpio_dm2[23]
port 324 nsew signal output
rlabel metal3 s -400 917228 60 917298 4 gpio_dm2[24]
port 325 nsew signal output
rlabel metal3 s -400 747428 60 747498 4 gpio_dm2[25]
port 326 nsew signal output
rlabel metal3 s -400 704228 60 704298 4 gpio_dm2[26]
port 327 nsew signal output
rlabel metal3 s -400 661028 60 661098 4 gpio_dm2[27]
port 328 nsew signal output
rlabel metal3 s -400 617828 60 617898 4 gpio_dm2[28]
port 329 nsew signal output
rlabel metal3 s -400 574628 60 574698 4 gpio_dm2[29]
port 330 nsew signal output
rlabel metal3 s 633266 158828 633726 158898 6 gpio_dm2[2]
port 331 nsew signal output
rlabel metal3 s -400 531428 60 531498 4 gpio_dm2[30]
port 332 nsew signal output
rlabel metal3 s -400 488228 60 488298 4 gpio_dm2[31]
port 333 nsew signal output
rlabel metal3 s -400 360628 60 360698 4 gpio_dm2[32]
port 334 nsew signal output
rlabel metal3 s -400 317428 60 317498 4 gpio_dm2[33]
port 335 nsew signal output
rlabel metal3 s -400 274228 60 274298 4 gpio_dm2[34]
port 336 nsew signal output
rlabel metal3 s -400 231028 60 231098 4 gpio_dm2[35]
port 337 nsew signal output
rlabel metal3 s -400 187828 60 187898 4 gpio_dm2[36]
port 338 nsew signal output
rlabel metal3 s -400 144628 60 144698 4 gpio_dm2[37]
port 339 nsew signal output
rlabel metal2 s 155034 -400 155090 56 8 gpio_dm2[38]
port 340 nsew signal output
rlabel metal2 s 263634 -400 263690 56 8 gpio_dm2[39]
port 341 nsew signal output
rlabel metal3 s 633266 204028 633726 204098 6 gpio_dm2[3]
port 342 nsew signal output
rlabel metal2 s 318434 -400 318490 56 8 gpio_dm2[40]
port 343 nsew signal output
rlabel metal2 s 373234 -400 373290 56 8 gpio_dm2[41]
port 344 nsew signal output
rlabel metal2 s 428034 -400 428090 56 8 gpio_dm2[42]
port 345 nsew signal output
rlabel metal2 s 482834 -400 482890 56 8 gpio_dm2[43]
port 346 nsew signal output
rlabel metal3 s 633266 249028 633726 249098 6 gpio_dm2[4]
port 347 nsew signal output
rlabel metal3 s 633266 294028 633726 294098 6 gpio_dm2[5]
port 348 nsew signal output
rlabel metal3 s 633266 339228 633726 339298 6 gpio_dm2[6]
port 349 nsew signal output
rlabel metal3 s 633266 516428 633726 516498 6 gpio_dm2[7]
port 350 nsew signal output
rlabel metal3 s 633266 561628 633726 561698 6 gpio_dm2[8]
port 351 nsew signal output
rlabel metal3 s 633266 606628 633726 606698 6 gpio_dm2[9]
port 352 nsew signal output
rlabel metal3 s 633266 69272 633726 69342 6 gpio_holdover[0]
port 353 nsew signal output
rlabel metal3 s 633266 652472 633726 652542 6 gpio_holdover[10]
port 354 nsew signal output
rlabel metal3 s 633266 697472 633726 697542 6 gpio_holdover[11]
port 355 nsew signal output
rlabel metal3 s 633266 742472 633726 742542 6 gpio_holdover[12]
port 356 nsew signal output
rlabel metal3 s 633206 831672 633726 831742 6 gpio_holdover[13]
port 357 nsew signal output
rlabel metal3 s 633266 920872 633726 920942 6 gpio_holdover[14]
port 358 nsew signal output
rlabel metal2 s 588392 953270 588448 953726 6 gpio_holdover[15]
port 359 nsew signal output
rlabel metal2 s 486592 953270 486648 953726 6 gpio_holdover[16]
port 360 nsew signal output
rlabel metal2 s 435192 953270 435248 953726 6 gpio_holdover[17]
port 361 nsew signal output
rlabel metal2 s 346192 953270 346248 953726 6 gpio_holdover[18]
port 362 nsew signal output
rlabel metal2 s 244392 953244 244448 953726 6 gpio_holdover[19]
port 363 nsew signal output
rlabel metal3 s 633266 114472 633726 114542 6 gpio_holdover[1]
port 364 nsew signal output
rlabel metal2 s 192792 953270 192848 953726 6 gpio_holdover[20]
port 365 nsew signal output
rlabel metal2 s 141392 953270 141448 953726 6 gpio_holdover[21]
port 366 nsew signal output
rlabel metal2 s 89992 953270 90048 953726 6 gpio_holdover[22]
port 367 nsew signal output
rlabel metal2 s 38592 953270 38648 953726 6 gpio_holdover[23]
port 368 nsew signal output
rlabel metal3 s -400 916584 60 916654 4 gpio_holdover[24]
port 369 nsew signal output
rlabel metal3 s -400 746784 60 746854 4 gpio_holdover[25]
port 370 nsew signal output
rlabel metal3 s -400 703584 60 703654 4 gpio_holdover[26]
port 371 nsew signal output
rlabel metal3 s -400 660384 60 660454 4 gpio_holdover[27]
port 372 nsew signal output
rlabel metal3 s -400 617184 60 617254 4 gpio_holdover[28]
port 373 nsew signal output
rlabel metal3 s -400 573984 60 574054 4 gpio_holdover[29]
port 374 nsew signal output
rlabel metal3 s 633266 159472 633726 159542 6 gpio_holdover[2]
port 375 nsew signal output
rlabel metal3 s -400 530784 60 530854 4 gpio_holdover[30]
port 376 nsew signal output
rlabel metal3 s -400 487584 60 487654 4 gpio_holdover[31]
port 377 nsew signal output
rlabel metal3 s -400 359984 60 360054 4 gpio_holdover[32]
port 378 nsew signal output
rlabel metal3 s -400 316784 60 316854 4 gpio_holdover[33]
port 379 nsew signal output
rlabel metal3 s -400 273584 60 273654 4 gpio_holdover[34]
port 380 nsew signal output
rlabel metal3 s -400 230384 60 230454 4 gpio_holdover[35]
port 381 nsew signal output
rlabel metal3 s -400 187184 60 187254 4 gpio_holdover[36]
port 382 nsew signal output
rlabel metal3 s -400 143984 60 144054 4 gpio_holdover[37]
port 383 nsew signal output
rlabel metal2 s 155678 -400 155734 56 8 gpio_holdover[38]
port 384 nsew signal output
rlabel metal2 s 264278 -400 264334 56 8 gpio_holdover[39]
port 385 nsew signal output
rlabel metal3 s 633266 204672 633726 204742 6 gpio_holdover[3]
port 386 nsew signal output
rlabel metal2 s 319078 -400 319134 56 8 gpio_holdover[40]
port 387 nsew signal output
rlabel metal2 s 373878 -400 373934 56 8 gpio_holdover[41]
port 388 nsew signal output
rlabel metal2 s 428678 -400 428734 56 8 gpio_holdover[42]
port 389 nsew signal output
rlabel metal2 s 483478 -400 483534 56 8 gpio_holdover[43]
port 390 nsew signal output
rlabel metal3 s 633266 249672 633726 249742 6 gpio_holdover[4]
port 391 nsew signal output
rlabel metal3 s 633266 294672 633726 294742 6 gpio_holdover[5]
port 392 nsew signal output
rlabel metal3 s 633266 339872 633726 339942 6 gpio_holdover[6]
port 393 nsew signal output
rlabel metal3 s 633266 517072 633726 517142 6 gpio_holdover[7]
port 394 nsew signal output
rlabel metal3 s 633266 562272 633726 562342 6 gpio_holdover[8]
port 395 nsew signal output
rlabel metal3 s 633266 607272 633726 607342 6 gpio_holdover[9]
port 396 nsew signal output
rlabel metal3 s 633266 72308 633726 72378 6 gpio_ib_mode_sel[0]
port 397 nsew signal output
rlabel metal3 s 633266 655508 633726 655578 6 gpio_ib_mode_sel[10]
port 398 nsew signal output
rlabel metal3 s 633266 700508 633726 700578 6 gpio_ib_mode_sel[11]
port 399 nsew signal output
rlabel metal3 s 633266 745508 633726 745578 6 gpio_ib_mode_sel[12]
port 400 nsew signal output
rlabel metal3 s 633266 834708 633726 834778 6 gpio_ib_mode_sel[13]
port 401 nsew signal output
rlabel metal3 s 633266 923908 633726 923978 6 gpio_ib_mode_sel[14]
port 402 nsew signal output
rlabel metal2 s 585356 953270 585412 953726 6 gpio_ib_mode_sel[15]
port 403 nsew signal output
rlabel metal2 s 483556 953270 483612 953726 6 gpio_ib_mode_sel[16]
port 404 nsew signal output
rlabel metal2 s 432156 953270 432212 953726 6 gpio_ib_mode_sel[17]
port 405 nsew signal output
rlabel metal2 s 343156 953270 343212 953726 6 gpio_ib_mode_sel[18]
port 406 nsew signal output
rlabel metal2 s 241356 953270 241412 953726 6 gpio_ib_mode_sel[19]
port 407 nsew signal output
rlabel metal3 s 633266 117508 633726 117578 6 gpio_ib_mode_sel[1]
port 408 nsew signal output
rlabel metal2 s 189756 953270 189812 953726 6 gpio_ib_mode_sel[20]
port 409 nsew signal output
rlabel metal2 s 138356 953270 138412 953726 6 gpio_ib_mode_sel[21]
port 410 nsew signal output
rlabel metal2 s 86956 953270 87012 953726 6 gpio_ib_mode_sel[22]
port 411 nsew signal output
rlabel metal2 s 35556 953270 35612 953726 6 gpio_ib_mode_sel[23]
port 412 nsew signal output
rlabel metal3 s -400 913548 60 913618 4 gpio_ib_mode_sel[24]
port 413 nsew signal output
rlabel metal3 s -400 743748 60 743818 4 gpio_ib_mode_sel[25]
port 414 nsew signal output
rlabel metal3 s -400 700548 60 700618 4 gpio_ib_mode_sel[26]
port 415 nsew signal output
rlabel metal3 s -400 657348 60 657418 4 gpio_ib_mode_sel[27]
port 416 nsew signal output
rlabel metal3 s -400 614148 60 614218 4 gpio_ib_mode_sel[28]
port 417 nsew signal output
rlabel metal3 s -400 570948 60 571018 4 gpio_ib_mode_sel[29]
port 418 nsew signal output
rlabel metal3 s 633266 162508 633726 162578 6 gpio_ib_mode_sel[2]
port 419 nsew signal output
rlabel metal3 s -400 527748 60 527818 4 gpio_ib_mode_sel[30]
port 420 nsew signal output
rlabel metal3 s -400 484548 60 484618 4 gpio_ib_mode_sel[31]
port 421 nsew signal output
rlabel metal3 s -400 356948 60 357018 4 gpio_ib_mode_sel[32]
port 422 nsew signal output
rlabel metal3 s -400 313748 60 313818 4 gpio_ib_mode_sel[33]
port 423 nsew signal output
rlabel metal3 s -400 270548 60 270618 4 gpio_ib_mode_sel[34]
port 424 nsew signal output
rlabel metal3 s -400 227348 60 227418 4 gpio_ib_mode_sel[35]
port 425 nsew signal output
rlabel metal3 s -400 184148 60 184218 4 gpio_ib_mode_sel[36]
port 426 nsew signal output
rlabel metal3 s -400 140948 60 141018 4 gpio_ib_mode_sel[37]
port 427 nsew signal output
rlabel metal2 s 158714 -400 158770 56 8 gpio_ib_mode_sel[38]
port 428 nsew signal output
rlabel metal2 s 267314 -400 267370 56 8 gpio_ib_mode_sel[39]
port 429 nsew signal output
rlabel metal3 s 633266 207708 633726 207778 6 gpio_ib_mode_sel[3]
port 430 nsew signal output
rlabel metal2 s 322114 -400 322170 56 8 gpio_ib_mode_sel[40]
port 431 nsew signal output
rlabel metal2 s 376914 -400 376970 56 8 gpio_ib_mode_sel[41]
port 432 nsew signal output
rlabel metal2 s 431714 -400 431770 56 8 gpio_ib_mode_sel[42]
port 433 nsew signal output
rlabel metal2 s 486514 -400 486570 56 8 gpio_ib_mode_sel[43]
port 434 nsew signal output
rlabel metal3 s 633266 252708 633726 252778 6 gpio_ib_mode_sel[4]
port 435 nsew signal output
rlabel metal3 s 633266 297708 633726 297778 6 gpio_ib_mode_sel[5]
port 436 nsew signal output
rlabel metal3 s 633266 342908 633726 342978 6 gpio_ib_mode_sel[6]
port 437 nsew signal output
rlabel metal3 s 633266 520108 633726 520178 6 gpio_ib_mode_sel[7]
port 438 nsew signal output
rlabel metal3 s 633266 565308 633726 565378 6 gpio_ib_mode_sel[8]
port 439 nsew signal output
rlabel metal3 s 633266 610308 633726 610378 6 gpio_ib_mode_sel[9]
port 440 nsew signal output
rlabel metal3 s 633266 58784 633726 58854 6 gpio_in[0]
port 441 nsew signal input
rlabel metal3 s 633266 641984 633726 642054 6 gpio_in[10]
port 442 nsew signal input
rlabel metal3 s 633266 686984 633726 687054 6 gpio_in[11]
port 443 nsew signal input
rlabel metal3 s 633266 731984 633726 732054 6 gpio_in[12]
port 444 nsew signal input
rlabel metal3 s 633266 821184 633726 821254 6 gpio_in[13]
port 445 nsew signal input
rlabel metal3 s 633266 910384 633726 910454 6 gpio_in[14]
port 446 nsew signal input
rlabel metal2 s 598880 953270 598936 953726 6 gpio_in[15]
port 447 nsew signal input
rlabel metal2 s 497080 953270 497136 953726 6 gpio_in[16]
port 448 nsew signal input
rlabel metal2 s 445680 953270 445736 953726 6 gpio_in[17]
port 449 nsew signal input
rlabel metal2 s 356680 953270 356736 953726 6 gpio_in[18]
port 450 nsew signal input
rlabel metal2 s 254880 953270 254936 953726 6 gpio_in[19]
port 451 nsew signal input
rlabel metal3 s 633266 103984 633726 104054 6 gpio_in[1]
port 452 nsew signal input
rlabel metal2 s 203280 953270 203336 953726 6 gpio_in[20]
port 453 nsew signal input
rlabel metal2 s 151880 953270 151936 953726 6 gpio_in[21]
port 454 nsew signal input
rlabel metal2 s 100480 953270 100536 953726 6 gpio_in[22]
port 455 nsew signal input
rlabel metal2 s 49080 953270 49136 953726 6 gpio_in[23]
port 456 nsew signal input
rlabel metal3 s -400 927072 60 927142 4 gpio_in[24]
port 457 nsew signal input
rlabel metal3 s -400 757272 60 757342 4 gpio_in[25]
port 458 nsew signal input
rlabel metal3 s -400 714072 60 714142 4 gpio_in[26]
port 459 nsew signal input
rlabel metal3 s -400 670872 60 670942 4 gpio_in[27]
port 460 nsew signal input
rlabel metal3 s -400 627672 60 627742 4 gpio_in[28]
port 461 nsew signal input
rlabel metal3 s -400 584472 60 584542 4 gpio_in[29]
port 462 nsew signal input
rlabel metal3 s 633266 148984 633726 149054 6 gpio_in[2]
port 463 nsew signal input
rlabel metal3 s -400 541272 60 541342 4 gpio_in[30]
port 464 nsew signal input
rlabel metal3 s -400 498072 60 498142 4 gpio_in[31]
port 465 nsew signal input
rlabel metal3 s -400 370472 60 370542 4 gpio_in[32]
port 466 nsew signal input
rlabel metal3 s -400 327272 60 327342 4 gpio_in[33]
port 467 nsew signal input
rlabel metal3 s -400 284072 60 284142 4 gpio_in[34]
port 468 nsew signal input
rlabel metal3 s -400 240872 60 240942 4 gpio_in[35]
port 469 nsew signal input
rlabel metal3 s -400 197672 60 197742 4 gpio_in[36]
port 470 nsew signal input
rlabel metal3 s -400 154472 60 154542 4 gpio_in[37]
port 471 nsew signal input
rlabel metal2 s 145190 -400 145246 56 8 gpio_in[38]
port 472 nsew signal input
rlabel metal2 s 253790 -400 253846 56 8 gpio_in[39]
port 473 nsew signal input
rlabel metal3 s 633266 194184 633726 194254 6 gpio_in[3]
port 474 nsew signal input
rlabel metal2 s 308590 -400 308646 56 8 gpio_in[40]
port 475 nsew signal input
rlabel metal2 s 363390 -400 363446 56 8 gpio_in[41]
port 476 nsew signal input
rlabel metal2 s 418190 -400 418246 56 8 gpio_in[42]
port 477 nsew signal input
rlabel metal2 s 472990 -400 473046 56 8 gpio_in[43]
port 478 nsew signal input
rlabel metal3 s 633266 239184 633726 239254 6 gpio_in[4]
port 479 nsew signal input
rlabel metal3 s 633266 284184 633726 284254 6 gpio_in[5]
port 480 nsew signal input
rlabel metal3 s 633266 329384 633726 329454 6 gpio_in[6]
port 481 nsew signal input
rlabel metal3 s 633266 506584 633726 506654 6 gpio_in[7]
port 482 nsew signal input
rlabel metal3 s 633266 551784 633726 551854 6 gpio_in[8]
port 483 nsew signal input
rlabel metal3 s 633266 596784 633726 596854 6 gpio_in[9]
port 484 nsew signal input
rlabel metal3 s 633266 73504 633726 73574 6 gpio_in_h[0]
port 485 nsew signal input
rlabel metal3 s 633266 656704 633726 656774 6 gpio_in_h[10]
port 486 nsew signal input
rlabel metal3 s 633266 701704 633726 701774 6 gpio_in_h[11]
port 487 nsew signal input
rlabel metal3 s 633266 746704 633726 746774 6 gpio_in_h[12]
port 488 nsew signal input
rlabel metal3 s 633266 835904 633726 835974 6 gpio_in_h[13]
port 489 nsew signal input
rlabel metal3 s 633266 925104 633726 925174 6 gpio_in_h[14]
port 490 nsew signal input
rlabel metal2 s 584160 953270 584216 953726 6 gpio_in_h[15]
port 491 nsew signal input
rlabel metal2 s 482360 953270 482416 953726 6 gpio_in_h[16]
port 492 nsew signal input
rlabel metal2 s 430960 953270 431016 953726 6 gpio_in_h[17]
port 493 nsew signal input
rlabel metal2 s 341960 953270 342016 953726 6 gpio_in_h[18]
port 494 nsew signal input
rlabel metal2 s 240160 953270 240216 953726 6 gpio_in_h[19]
port 495 nsew signal input
rlabel metal3 s 633266 118704 633726 118774 6 gpio_in_h[1]
port 496 nsew signal input
rlabel metal2 s 188560 953270 188616 953726 6 gpio_in_h[20]
port 497 nsew signal input
rlabel metal2 s 137160 953270 137216 953726 6 gpio_in_h[21]
port 498 nsew signal input
rlabel metal2 s 85760 953270 85816 953726 6 gpio_in_h[22]
port 499 nsew signal input
rlabel metal2 s 34360 953270 34416 953726 6 gpio_in_h[23]
port 500 nsew signal input
rlabel metal3 s -400 912352 60 912422 4 gpio_in_h[24]
port 501 nsew signal input
rlabel metal3 s -400 742552 60 742622 4 gpio_in_h[25]
port 502 nsew signal input
rlabel metal3 s -400 699352 60 699422 4 gpio_in_h[26]
port 503 nsew signal input
rlabel metal3 s -400 656152 60 656222 4 gpio_in_h[27]
port 504 nsew signal input
rlabel metal3 s -400 612952 60 613022 4 gpio_in_h[28]
port 505 nsew signal input
rlabel metal3 s -400 569752 60 569822 4 gpio_in_h[29]
port 506 nsew signal input
rlabel metal3 s 633266 163704 633726 163774 6 gpio_in_h[2]
port 507 nsew signal input
rlabel metal3 s -400 526552 60 526622 4 gpio_in_h[30]
port 508 nsew signal input
rlabel metal3 s -400 483352 60 483422 4 gpio_in_h[31]
port 509 nsew signal input
rlabel metal3 s -400 355752 60 355822 4 gpio_in_h[32]
port 510 nsew signal input
rlabel metal3 s -400 312552 60 312622 4 gpio_in_h[33]
port 511 nsew signal input
rlabel metal3 s -400 269352 60 269422 4 gpio_in_h[34]
port 512 nsew signal input
rlabel metal3 s -400 226152 60 226222 4 gpio_in_h[35]
port 513 nsew signal input
rlabel metal3 s -400 182952 60 183022 4 gpio_in_h[36]
port 514 nsew signal input
rlabel metal3 s -400 139752 60 139822 4 gpio_in_h[37]
port 515 nsew signal input
rlabel metal2 s 159910 -400 159966 56 8 gpio_in_h[38]
port 516 nsew signal input
rlabel metal2 s 268510 -400 268566 56 8 gpio_in_h[39]
port 517 nsew signal input
rlabel metal3 s 633266 208904 633726 208974 6 gpio_in_h[3]
port 518 nsew signal input
rlabel metal2 s 323310 -400 323366 56 8 gpio_in_h[40]
port 519 nsew signal input
rlabel metal2 s 378110 -400 378166 56 8 gpio_in_h[41]
port 520 nsew signal input
rlabel metal2 s 432910 -400 432966 56 8 gpio_in_h[42]
port 521 nsew signal input
rlabel metal2 s 487710 -400 487766 56 8 gpio_in_h[43]
port 522 nsew signal input
rlabel metal3 s 633266 253904 633726 253974 6 gpio_in_h[4]
port 523 nsew signal input
rlabel metal3 s 633266 298904 633726 298974 6 gpio_in_h[5]
port 524 nsew signal input
rlabel metal3 s 633266 344104 633726 344174 6 gpio_in_h[6]
port 525 nsew signal input
rlabel metal3 s 633266 521304 633726 521374 6 gpio_in_h[7]
port 526 nsew signal input
rlabel metal3 s 633266 566504 633726 566574 6 gpio_in_h[8]
port 527 nsew signal input
rlabel metal3 s 633266 611504 633726 611574 6 gpio_in_h[9]
port 528 nsew signal input
rlabel metal3 s 633266 65500 633726 65570 6 gpio_inp_dis[0]
port 529 nsew signal output
rlabel metal3 s 633266 648700 633726 648770 6 gpio_inp_dis[10]
port 530 nsew signal output
rlabel metal3 s 633266 693700 633726 693770 6 gpio_inp_dis[11]
port 531 nsew signal output
rlabel metal3 s 633266 738700 633726 738770 6 gpio_inp_dis[12]
port 532 nsew signal output
rlabel metal3 s 633266 827900 633726 827970 6 gpio_inp_dis[13]
port 533 nsew signal output
rlabel metal3 s 633266 917100 633726 917170 6 gpio_inp_dis[14]
port 534 nsew signal output
rlabel metal2 s 592164 953270 592220 953726 6 gpio_inp_dis[15]
port 535 nsew signal output
rlabel metal2 s 490364 953270 490420 953726 6 gpio_inp_dis[16]
port 536 nsew signal output
rlabel metal2 s 438964 953270 439020 953726 6 gpio_inp_dis[17]
port 537 nsew signal output
rlabel metal2 s 349964 953270 350020 953726 6 gpio_inp_dis[18]
port 538 nsew signal output
rlabel metal2 s 248164 953270 248220 953726 6 gpio_inp_dis[19]
port 539 nsew signal output
rlabel metal3 s 633266 110700 633726 110770 6 gpio_inp_dis[1]
port 540 nsew signal output
rlabel metal2 s 196564 953270 196620 953726 6 gpio_inp_dis[20]
port 541 nsew signal output
rlabel metal2 s 145164 953270 145220 953726 6 gpio_inp_dis[21]
port 542 nsew signal output
rlabel metal2 s 93764 953270 93820 953726 6 gpio_inp_dis[22]
port 543 nsew signal output
rlabel metal2 s 42364 953270 42420 953726 6 gpio_inp_dis[23]
port 544 nsew signal output
rlabel metal3 s -400 920356 60 920426 4 gpio_inp_dis[24]
port 545 nsew signal output
rlabel metal3 s -400 750556 60 750626 4 gpio_inp_dis[25]
port 546 nsew signal output
rlabel metal3 s -400 707356 60 707426 4 gpio_inp_dis[26]
port 547 nsew signal output
rlabel metal3 s -400 664156 60 664226 4 gpio_inp_dis[27]
port 548 nsew signal output
rlabel metal3 s -400 620956 60 621026 4 gpio_inp_dis[28]
port 549 nsew signal output
rlabel metal3 s -400 577756 60 577826 4 gpio_inp_dis[29]
port 550 nsew signal output
rlabel metal3 s 633266 155700 633726 155770 6 gpio_inp_dis[2]
port 551 nsew signal output
rlabel metal3 s -400 534556 60 534626 4 gpio_inp_dis[30]
port 552 nsew signal output
rlabel metal3 s -400 491356 60 491426 4 gpio_inp_dis[31]
port 553 nsew signal output
rlabel metal3 s -400 363756 60 363826 4 gpio_inp_dis[32]
port 554 nsew signal output
rlabel metal3 s -400 320556 60 320626 4 gpio_inp_dis[33]
port 555 nsew signal output
rlabel metal3 s -400 277356 60 277426 4 gpio_inp_dis[34]
port 556 nsew signal output
rlabel metal3 s -400 234156 60 234226 4 gpio_inp_dis[35]
port 557 nsew signal output
rlabel metal3 s -400 190956 60 191026 4 gpio_inp_dis[36]
port 558 nsew signal output
rlabel metal3 s -400 147756 60 147826 4 gpio_inp_dis[37]
port 559 nsew signal output
rlabel metal2 s 151906 -400 151962 56 8 gpio_inp_dis[38]
port 560 nsew signal output
rlabel metal2 s 260506 -400 260562 56 8 gpio_inp_dis[39]
port 561 nsew signal output
rlabel metal3 s 633266 200900 633726 200970 6 gpio_inp_dis[3]
port 562 nsew signal output
rlabel metal2 s 315306 -400 315362 56 8 gpio_inp_dis[40]
port 563 nsew signal output
rlabel metal2 s 370106 -400 370162 56 8 gpio_inp_dis[41]
port 564 nsew signal output
rlabel metal2 s 424906 -400 424962 56 8 gpio_inp_dis[42]
port 565 nsew signal output
rlabel metal2 s 479706 -400 479762 56 8 gpio_inp_dis[43]
port 566 nsew signal output
rlabel metal3 s 633266 245900 633726 245970 6 gpio_inp_dis[4]
port 567 nsew signal output
rlabel metal3 s 633266 290900 633726 290970 6 gpio_inp_dis[5]
port 568 nsew signal output
rlabel metal3 s 633266 336100 633726 336170 6 gpio_inp_dis[6]
port 569 nsew signal output
rlabel metal3 s 633266 513300 633726 513370 6 gpio_inp_dis[7]
port 570 nsew signal output
rlabel metal3 s 633266 558500 633726 558570 6 gpio_inp_dis[8]
port 571 nsew signal output
rlabel metal3 s 633266 603500 633726 603570 6 gpio_inp_dis[9]
port 572 nsew signal output
rlabel metal3 s 633266 76005 633726 76067 6 gpio_loopback_one[0]
port 573 nsew signal input
rlabel metal3 s 633266 658006 633726 658068 6 gpio_loopback_one[10]
port 574 nsew signal input
rlabel metal3 s 633266 703006 633726 703068 6 gpio_loopback_one[11]
port 575 nsew signal input
rlabel metal3 s 633266 748006 633726 748068 6 gpio_loopback_one[12]
port 576 nsew signal input
rlabel metal3 s 633266 837006 633726 837068 6 gpio_loopback_one[13]
port 577 nsew signal input
rlabel metal3 s 633266 927006 633726 927068 6 gpio_loopback_one[14]
port 578 nsew signal input
rlabel metal2 s 578298 953270 578358 953726 6 gpio_loopback_one[15]
port 579 nsew signal input
rlabel metal2 s 478898 953270 478958 953726 6 gpio_loopback_one[16]
port 580 nsew signal input
rlabel metal2 s 427698 953270 427758 953726 6 gpio_loopback_one[17]
port 581 nsew signal input
rlabel metal2 s 338698 953270 338758 953726 6 gpio_loopback_one[18]
port 582 nsew signal input
rlabel metal2 s 234298 953270 234358 953726 6 gpio_loopback_one[19]
port 583 nsew signal input
rlabel metal3 s 633266 121005 633726 121067 6 gpio_loopback_one[1]
port 584 nsew signal input
rlabel metal2 s 183098 953270 183158 953726 6 gpio_loopback_one[20]
port 585 nsew signal input
rlabel metal2 s 131898 953270 131958 953726 6 gpio_loopback_one[21]
port 586 nsew signal input
rlabel metal2 s 80698 953270 80758 953726 6 gpio_loopback_one[22]
port 587 nsew signal input
rlabel metal2 s 29498 953270 29558 953726 6 gpio_loopback_one[23]
port 588 nsew signal input
rlabel metal3 s -400 906644 60 906704 4 gpio_loopback_one[24]
port 589 nsew signal input
rlabel metal3 s -400 736644 60 736704 4 gpio_loopback_one[25]
port 590 nsew signal input
rlabel metal3 s -400 693644 60 693704 4 gpio_loopback_one[26]
port 591 nsew signal input
rlabel metal3 s -400 650644 60 650704 4 gpio_loopback_one[27]
port 592 nsew signal input
rlabel metal3 s -400 607644 60 607704 4 gpio_loopback_one[28]
port 593 nsew signal input
rlabel metal3 s -400 564644 60 564704 4 gpio_loopback_one[29]
port 594 nsew signal input
rlabel metal3 s 633266 166005 633726 166067 6 gpio_loopback_one[2]
port 595 nsew signal input
rlabel metal3 s -400 521644 60 521704 4 gpio_loopback_one[30]
port 596 nsew signal input
rlabel metal3 s -400 478644 60 478704 4 gpio_loopback_one[31]
port 597 nsew signal input
rlabel metal3 s -400 349644 60 349704 4 gpio_loopback_one[32]
port 598 nsew signal input
rlabel metal3 s -400 306644 60 306704 4 gpio_loopback_one[33]
port 599 nsew signal input
rlabel metal3 s -400 263644 60 263704 4 gpio_loopback_one[34]
port 600 nsew signal input
rlabel metal3 s -400 220644 60 220704 4 gpio_loopback_one[35]
port 601 nsew signal input
rlabel metal3 s -400 177644 60 177704 4 gpio_loopback_one[36]
port 602 nsew signal input
rlabel metal3 s -400 134644 60 134704 4 gpio_loopback_one[37]
port 603 nsew signal input
rlabel metal2 s 160580 -400 160632 56 8 gpio_loopback_one[38]
port 604 nsew signal input
rlabel metal2 s 269180 -400 269232 56 8 gpio_loopback_one[39]
port 605 nsew signal input
rlabel metal3 s 633266 211005 633726 211067 6 gpio_loopback_one[3]
port 606 nsew signal input
rlabel metal2 s 323980 -400 324032 56 8 gpio_loopback_one[40]
port 607 nsew signal input
rlabel metal2 s 378780 -400 378832 56 8 gpio_loopback_one[41]
port 608 nsew signal input
rlabel metal2 s 433580 -400 433632 56 8 gpio_loopback_one[42]
port 609 nsew signal input
rlabel metal2 s 488380 -400 488432 56 8 gpio_loopback_one[43]
port 610 nsew signal input
rlabel metal3 s 633266 256005 633726 256067 6 gpio_loopback_one[4]
port 611 nsew signal input
rlabel metal3 s 633266 301005 633726 301067 6 gpio_loopback_one[5]
port 612 nsew signal input
rlabel metal3 s 633266 346005 633726 346067 6 gpio_loopback_one[6]
port 613 nsew signal input
rlabel metal3 s 633266 523005 633726 523067 6 gpio_loopback_one[7]
port 614 nsew signal input
rlabel metal3 s 633266 568006 633726 568068 6 gpio_loopback_one[8]
port 615 nsew signal input
rlabel metal3 s 633266 613006 633726 613068 6 gpio_loopback_one[9]
port 616 nsew signal input
rlabel metal3 s 633266 78006 633726 78068 6 gpio_loopback_zero[0]
port 617 nsew signal input
rlabel metal3 s 633266 660006 633726 660068 6 gpio_loopback_zero[10]
port 618 nsew signal input
rlabel metal3 s 633266 705006 633726 705068 6 gpio_loopback_zero[11]
port 619 nsew signal input
rlabel metal3 s 633266 750006 633726 750068 6 gpio_loopback_zero[12]
port 620 nsew signal input
rlabel metal3 s 633266 839006 633726 839068 6 gpio_loopback_zero[13]
port 621 nsew signal input
rlabel metal3 s 633266 929006 633726 929068 6 gpio_loopback_zero[14]
port 622 nsew signal input
rlabel metal2 s 576298 953270 576358 953726 6 gpio_loopback_zero[15]
port 623 nsew signal input
rlabel metal2 s 476898 953270 476958 953726 6 gpio_loopback_zero[16]
port 624 nsew signal input
rlabel metal2 s 425698 953270 425758 953726 6 gpio_loopback_zero[17]
port 625 nsew signal input
rlabel metal2 s 336698 953270 336758 953726 6 gpio_loopback_zero[18]
port 626 nsew signal input
rlabel metal2 s 232298 953270 232358 953726 6 gpio_loopback_zero[19]
port 627 nsew signal input
rlabel metal3 s 633266 123006 633726 123068 6 gpio_loopback_zero[1]
port 628 nsew signal input
rlabel metal2 s 181098 953270 181158 953726 6 gpio_loopback_zero[20]
port 629 nsew signal input
rlabel metal2 s 129898 953270 129958 953726 6 gpio_loopback_zero[21]
port 630 nsew signal input
rlabel metal2 s 78698 953270 78758 953726 6 gpio_loopback_zero[22]
port 631 nsew signal input
rlabel metal2 s 27498 953270 27558 953726 6 gpio_loopback_zero[23]
port 632 nsew signal input
rlabel metal3 s -400 904644 122 904704 4 gpio_loopback_zero[24]
port 633 nsew signal input
rlabel metal3 s -400 734644 122 734704 4 gpio_loopback_zero[25]
port 634 nsew signal input
rlabel metal3 s -400 691644 674 691704 6 gpio_loopback_zero[26]
port 635 nsew signal input
rlabel metal3 s -400 648644 674 648704 6 gpio_loopback_zero[27]
port 636 nsew signal input
rlabel metal3 s -400 605644 674 605704 6 gpio_loopback_zero[28]
port 637 nsew signal input
rlabel metal3 s -400 562644 674 562704 6 gpio_loopback_zero[29]
port 638 nsew signal input
rlabel metal3 s 633266 168006 633726 168068 6 gpio_loopback_zero[2]
port 639 nsew signal input
rlabel metal3 s -400 519644 674 519704 6 gpio_loopback_zero[30]
port 640 nsew signal input
rlabel metal3 s -400 476644 674 476704 6 gpio_loopback_zero[31]
port 641 nsew signal input
rlabel metal3 s -400 347644 674 347704 6 gpio_loopback_zero[32]
port 642 nsew signal input
rlabel metal3 s -400 304644 674 304704 6 gpio_loopback_zero[33]
port 643 nsew signal input
rlabel metal3 s -400 261644 674 261704 6 gpio_loopback_zero[34]
port 644 nsew signal input
rlabel metal3 s -400 218644 674 218704 6 gpio_loopback_zero[35]
port 645 nsew signal input
rlabel metal3 s -400 175644 674 175704 6 gpio_loopback_zero[36]
port 646 nsew signal input
rlabel metal3 s -400 132644 674 132704 6 gpio_loopback_zero[37]
port 647 nsew signal input
rlabel metal2 s 163791 -400 163843 56 8 gpio_loopback_zero[38]
port 648 nsew signal input
rlabel metal2 s 273360 -400 273412 56 8 gpio_loopback_zero[39]
port 649 nsew signal input
rlabel metal3 s 633266 213006 633726 213068 6 gpio_loopback_zero[3]
port 650 nsew signal input
rlabel metal2 s 328165 -400 328217 56 8 gpio_loopback_zero[40]
port 651 nsew signal input
rlabel metal2 s 382978 -400 383030 56 8 gpio_loopback_zero[41]
port 652 nsew signal input
rlabel metal2 s 437778 -400 437830 56 8 gpio_loopback_zero[42]
port 653 nsew signal input
rlabel metal2 s 492635 -400 492687 56 8 gpio_loopback_zero[43]
port 654 nsew signal input
rlabel metal3 s 633266 258006 633726 258068 6 gpio_loopback_zero[4]
port 655 nsew signal input
rlabel metal3 s 633266 303006 633726 303068 6 gpio_loopback_zero[5]
port 656 nsew signal input
rlabel metal3 s 633266 348006 633726 348068 6 gpio_loopback_zero[6]
port 657 nsew signal input
rlabel metal3 s 633266 525006 633726 525068 6 gpio_loopback_zero[7]
port 658 nsew signal input
rlabel metal3 s 633266 570006 633726 570068 6 gpio_loopback_zero[8]
port 659 nsew signal input
rlabel metal3 s 633266 615006 633726 615068 6 gpio_loopback_zero[9]
port 660 nsew signal input
rlabel metal3 s 633266 72952 633726 73022 6 gpio_oeb[0]
port 661 nsew signal output
rlabel metal3 s 633266 656152 633726 656222 6 gpio_oeb[10]
port 662 nsew signal output
rlabel metal3 s 633266 701152 633726 701222 6 gpio_oeb[11]
port 663 nsew signal output
rlabel metal3 s 633266 746152 633726 746222 6 gpio_oeb[12]
port 664 nsew signal output
rlabel metal3 s 633266 835352 633726 835422 6 gpio_oeb[13]
port 665 nsew signal output
rlabel metal3 s 633266 924552 633726 924622 6 gpio_oeb[14]
port 666 nsew signal output
rlabel metal2 s 584712 953270 584768 953726 6 gpio_oeb[15]
port 667 nsew signal output
rlabel metal2 s 482912 953270 482968 953726 6 gpio_oeb[16]
port 668 nsew signal output
rlabel metal2 s 431512 953270 431568 953726 6 gpio_oeb[17]
port 669 nsew signal output
rlabel metal2 s 342512 953270 342568 953726 6 gpio_oeb[18]
port 670 nsew signal output
rlabel metal2 s 240712 953270 240768 953726 6 gpio_oeb[19]
port 671 nsew signal output
rlabel metal3 s 633266 118152 633726 118222 6 gpio_oeb[1]
port 672 nsew signal output
rlabel metal2 s 189112 953270 189168 953726 6 gpio_oeb[20]
port 673 nsew signal output
rlabel metal2 s 137712 953270 137768 953726 6 gpio_oeb[21]
port 674 nsew signal output
rlabel metal2 s 86312 953270 86368 953726 6 gpio_oeb[22]
port 675 nsew signal output
rlabel metal2 s 34912 953270 34968 953726 6 gpio_oeb[23]
port 676 nsew signal output
rlabel metal3 s -400 912904 60 912974 4 gpio_oeb[24]
port 677 nsew signal output
rlabel metal3 s -400 743104 60 743174 4 gpio_oeb[25]
port 678 nsew signal output
rlabel metal3 s -400 699904 60 699974 4 gpio_oeb[26]
port 679 nsew signal output
rlabel metal3 s -400 656704 60 656774 4 gpio_oeb[27]
port 680 nsew signal output
rlabel metal3 s -400 613504 60 613574 4 gpio_oeb[28]
port 681 nsew signal output
rlabel metal3 s -400 570304 60 570374 4 gpio_oeb[29]
port 682 nsew signal output
rlabel metal3 s 633266 163152 633726 163222 6 gpio_oeb[2]
port 683 nsew signal output
rlabel metal3 s -400 527104 60 527174 4 gpio_oeb[30]
port 684 nsew signal output
rlabel metal3 s -400 483904 60 483974 4 gpio_oeb[31]
port 685 nsew signal output
rlabel metal3 s -400 356304 60 356374 4 gpio_oeb[32]
port 686 nsew signal output
rlabel metal3 s -400 313104 60 313174 4 gpio_oeb[33]
port 687 nsew signal output
rlabel metal3 s -400 269904 60 269974 4 gpio_oeb[34]
port 688 nsew signal output
rlabel metal3 s -400 226704 60 226774 4 gpio_oeb[35]
port 689 nsew signal output
rlabel metal3 s -400 183504 60 183574 4 gpio_oeb[36]
port 690 nsew signal output
rlabel metal3 s -400 140304 60 140374 4 gpio_oeb[37]
port 691 nsew signal output
rlabel metal2 s 159358 -400 159414 56 8 gpio_oeb[38]
port 692 nsew signal output
rlabel metal2 s 267958 -400 268014 56 8 gpio_oeb[39]
port 693 nsew signal output
rlabel metal3 s 633266 208352 633726 208422 6 gpio_oeb[3]
port 694 nsew signal output
rlabel metal2 s 322758 -400 322814 56 8 gpio_oeb[40]
port 695 nsew signal output
rlabel metal2 s 377558 -400 377614 56 8 gpio_oeb[41]
port 696 nsew signal output
rlabel metal2 s 432358 -400 432414 56 8 gpio_oeb[42]
port 697 nsew signal output
rlabel metal2 s 487158 -400 487214 56 8 gpio_oeb[43]
port 698 nsew signal output
rlabel metal3 s 633266 253352 633726 253422 6 gpio_oeb[4]
port 699 nsew signal output
rlabel metal3 s 633266 298352 633726 298422 6 gpio_oeb[5]
port 700 nsew signal output
rlabel metal3 s 633266 343552 633726 343622 6 gpio_oeb[6]
port 701 nsew signal output
rlabel metal3 s 633266 520752 633726 520822 6 gpio_oeb[7]
port 702 nsew signal output
rlabel metal3 s 633266 565952 633726 566022 6 gpio_oeb[8]
port 703 nsew signal output
rlabel metal3 s 633266 610952 633726 611022 6 gpio_oeb[9]
port 704 nsew signal output
rlabel metal3 s 633266 69824 633726 69894 6 gpio_out[0]
port 705 nsew signal output
rlabel metal3 s 633266 653024 633726 653094 6 gpio_out[10]
port 706 nsew signal output
rlabel metal3 s 633266 698024 633726 698094 6 gpio_out[11]
port 707 nsew signal output
rlabel metal3 s 633266 743024 633726 743094 6 gpio_out[12]
port 708 nsew signal output
rlabel metal3 s 633266 832224 633726 832294 6 gpio_out[13]
port 709 nsew signal output
rlabel metal3 s 633266 921424 633726 921494 6 gpio_out[14]
port 710 nsew signal output
rlabel metal2 s 587840 953270 587896 953726 6 gpio_out[15]
port 711 nsew signal output
rlabel metal2 s 486040 953270 486096 953726 6 gpio_out[16]
port 712 nsew signal output
rlabel metal2 s 434640 953270 434696 953726 6 gpio_out[17]
port 713 nsew signal output
rlabel metal2 s 345640 953270 345696 953726 6 gpio_out[18]
port 714 nsew signal output
rlabel metal2 s 243840 953270 243896 953726 6 gpio_out[19]
port 715 nsew signal output
rlabel metal3 s 633266 115024 633726 115094 6 gpio_out[1]
port 716 nsew signal output
rlabel metal2 s 192240 953270 192296 953726 6 gpio_out[20]
port 717 nsew signal output
rlabel metal2 s 140840 953270 140896 953726 6 gpio_out[21]
port 718 nsew signal output
rlabel metal2 s 89440 953270 89496 953726 6 gpio_out[22]
port 719 nsew signal output
rlabel metal2 s 38040 953270 38096 953726 6 gpio_out[23]
port 720 nsew signal output
rlabel metal3 s -400 916032 60 916102 4 gpio_out[24]
port 721 nsew signal output
rlabel metal3 s -400 746232 60 746302 4 gpio_out[25]
port 722 nsew signal output
rlabel metal3 s -400 703032 60 703102 4 gpio_out[26]
port 723 nsew signal output
rlabel metal3 s -400 659832 60 659902 4 gpio_out[27]
port 724 nsew signal output
rlabel metal3 s -400 616632 60 616702 4 gpio_out[28]
port 725 nsew signal output
rlabel metal3 s -400 573432 60 573502 4 gpio_out[29]
port 726 nsew signal output
rlabel metal3 s 633266 160024 633726 160094 6 gpio_out[2]
port 727 nsew signal output
rlabel metal3 s -400 530232 60 530302 4 gpio_out[30]
port 728 nsew signal output
rlabel metal3 s -400 487032 60 487102 4 gpio_out[31]
port 729 nsew signal output
rlabel metal3 s -400 359432 60 359502 4 gpio_out[32]
port 730 nsew signal output
rlabel metal3 s -400 316232 60 316302 4 gpio_out[33]
port 731 nsew signal output
rlabel metal3 s -400 273032 60 273102 4 gpio_out[34]
port 732 nsew signal output
rlabel metal3 s -400 229832 60 229902 4 gpio_out[35]
port 733 nsew signal output
rlabel metal3 s -400 186632 60 186702 4 gpio_out[36]
port 734 nsew signal output
rlabel metal3 s -400 143432 60 143502 4 gpio_out[37]
port 735 nsew signal output
rlabel metal2 s 156230 -400 156286 56 8 gpio_out[38]
port 736 nsew signal output
rlabel metal2 s 264830 -400 264886 56 8 gpio_out[39]
port 737 nsew signal output
rlabel metal3 s 633266 205224 633726 205294 6 gpio_out[3]
port 738 nsew signal output
rlabel metal2 s 319630 -400 319686 56 8 gpio_out[40]
port 739 nsew signal output
rlabel metal2 s 374430 -400 374486 56 8 gpio_out[41]
port 740 nsew signal output
rlabel metal2 s 429230 -400 429286 56 8 gpio_out[42]
port 741 nsew signal output
rlabel metal2 s 484030 -400 484086 56 8 gpio_out[43]
port 742 nsew signal output
rlabel metal3 s 633266 250224 633726 250294 6 gpio_out[4]
port 743 nsew signal output
rlabel metal3 s 633266 295224 633726 295294 6 gpio_out[5]
port 744 nsew signal output
rlabel metal3 s 633266 340424 633726 340494 6 gpio_out[6]
port 745 nsew signal output
rlabel metal3 s 633266 517624 633726 517694 6 gpio_out[7]
port 746 nsew signal output
rlabel metal3 s 633266 562824 633726 562894 6 gpio_out[8]
port 747 nsew signal output
rlabel metal3 s 633266 607824 633726 607894 6 gpio_out[9]
port 748 nsew signal output
rlabel metal3 s 633266 60624 633726 60694 6 gpio_slow_sel[0]
port 749 nsew signal output
rlabel metal3 s 633266 643824 633726 643894 6 gpio_slow_sel[10]
port 750 nsew signal output
rlabel metal3 s 633266 688824 633726 688894 6 gpio_slow_sel[11]
port 751 nsew signal output
rlabel metal3 s 633266 733824 633726 733894 6 gpio_slow_sel[12]
port 752 nsew signal output
rlabel metal3 s 633266 823024 633726 823094 6 gpio_slow_sel[13]
port 753 nsew signal output
rlabel metal3 s 633266 912224 633726 912294 6 gpio_slow_sel[14]
port 754 nsew signal output
rlabel metal2 s 597040 953270 597096 953726 6 gpio_slow_sel[15]
port 755 nsew signal output
rlabel metal2 s 495240 953270 495296 953726 6 gpio_slow_sel[16]
port 756 nsew signal output
rlabel metal2 s 443840 953270 443896 953726 6 gpio_slow_sel[17]
port 757 nsew signal output
rlabel metal2 s 354840 953270 354896 953726 6 gpio_slow_sel[18]
port 758 nsew signal output
rlabel metal2 s 253040 953270 253096 953726 6 gpio_slow_sel[19]
port 759 nsew signal output
rlabel metal3 s 633266 105824 633726 105894 6 gpio_slow_sel[1]
port 760 nsew signal output
rlabel metal2 s 201440 953270 201496 953726 6 gpio_slow_sel[20]
port 761 nsew signal output
rlabel metal2 s 150040 953270 150096 953726 6 gpio_slow_sel[21]
port 762 nsew signal output
rlabel metal2 s 98640 953270 98696 953726 6 gpio_slow_sel[22]
port 763 nsew signal output
rlabel metal2 s 47240 953270 47296 953726 6 gpio_slow_sel[23]
port 764 nsew signal output
rlabel metal3 s -400 925232 60 925302 4 gpio_slow_sel[24]
port 765 nsew signal output
rlabel metal3 s -400 755432 60 755502 4 gpio_slow_sel[25]
port 766 nsew signal output
rlabel metal3 s -400 712232 60 712302 4 gpio_slow_sel[26]
port 767 nsew signal output
rlabel metal3 s -400 669032 60 669102 4 gpio_slow_sel[27]
port 768 nsew signal output
rlabel metal3 s -400 625832 60 625902 4 gpio_slow_sel[28]
port 769 nsew signal output
rlabel metal3 s -400 582632 60 582702 4 gpio_slow_sel[29]
port 770 nsew signal output
rlabel metal3 s 633266 150824 633726 150894 6 gpio_slow_sel[2]
port 771 nsew signal output
rlabel metal3 s -400 539432 60 539502 4 gpio_slow_sel[30]
port 772 nsew signal output
rlabel metal3 s -400 496232 60 496302 4 gpio_slow_sel[31]
port 773 nsew signal output
rlabel metal3 s -400 368632 60 368702 4 gpio_slow_sel[32]
port 774 nsew signal output
rlabel metal3 s -400 325432 60 325502 4 gpio_slow_sel[33]
port 775 nsew signal output
rlabel metal3 s -400 282232 60 282302 4 gpio_slow_sel[34]
port 776 nsew signal output
rlabel metal3 s -400 239032 60 239102 4 gpio_slow_sel[35]
port 777 nsew signal output
rlabel metal3 s -400 195832 60 195902 4 gpio_slow_sel[36]
port 778 nsew signal output
rlabel metal3 s -400 152632 60 152702 4 gpio_slow_sel[37]
port 779 nsew signal output
rlabel metal2 s 147030 -400 147086 56 8 gpio_slow_sel[38]
port 780 nsew signal output
rlabel metal2 s 255630 -400 255686 56 8 gpio_slow_sel[39]
port 781 nsew signal output
rlabel metal3 s 633266 196024 633726 196094 6 gpio_slow_sel[3]
port 782 nsew signal output
rlabel metal2 s 310430 -400 310486 56 8 gpio_slow_sel[40]
port 783 nsew signal output
rlabel metal2 s 365230 -400 365286 56 8 gpio_slow_sel[41]
port 784 nsew signal output
rlabel metal2 s 420030 -400 420086 56 8 gpio_slow_sel[42]
port 785 nsew signal output
rlabel metal2 s 474830 -400 474886 56 8 gpio_slow_sel[43]
port 786 nsew signal output
rlabel metal3 s 633266 241024 633726 241094 6 gpio_slow_sel[4]
port 787 nsew signal output
rlabel metal3 s 633266 286024 633726 286094 6 gpio_slow_sel[5]
port 788 nsew signal output
rlabel metal3 s 633266 331224 633726 331294 6 gpio_slow_sel[6]
port 789 nsew signal output
rlabel metal3 s 633266 508424 633726 508494 6 gpio_slow_sel[7]
port 790 nsew signal output
rlabel metal3 s 633266 553624 633726 553694 6 gpio_slow_sel[8]
port 791 nsew signal output
rlabel metal3 s 633266 598624 633726 598694 6 gpio_slow_sel[9]
port 792 nsew signal output
rlabel metal3 s 633266 71664 633726 71734 6 gpio_vtrip_sel[0]
port 793 nsew signal output
rlabel metal3 s 633266 654864 633726 654934 6 gpio_vtrip_sel[10]
port 794 nsew signal output
rlabel metal3 s 633266 699864 633726 699934 6 gpio_vtrip_sel[11]
port 795 nsew signal output
rlabel metal3 s 633266 744864 633726 744934 6 gpio_vtrip_sel[12]
port 796 nsew signal output
rlabel metal3 s 633266 834064 633726 834134 6 gpio_vtrip_sel[13]
port 797 nsew signal output
rlabel metal3 s 633266 923264 633726 923334 6 gpio_vtrip_sel[14]
port 798 nsew signal output
rlabel metal2 s 586000 953270 586056 953726 6 gpio_vtrip_sel[15]
port 799 nsew signal output
rlabel metal2 s 484200 953270 484256 953726 6 gpio_vtrip_sel[16]
port 800 nsew signal output
rlabel metal2 s 432800 953270 432856 953726 6 gpio_vtrip_sel[17]
port 801 nsew signal output
rlabel metal2 s 343800 953270 343856 953726 6 gpio_vtrip_sel[18]
port 802 nsew signal output
rlabel metal2 s 242000 953270 242056 953726 6 gpio_vtrip_sel[19]
port 803 nsew signal output
rlabel metal3 s 633266 116864 633726 116934 6 gpio_vtrip_sel[1]
port 804 nsew signal output
rlabel metal2 s 190400 953270 190456 953726 6 gpio_vtrip_sel[20]
port 805 nsew signal output
rlabel metal2 s 139000 953270 139056 953726 6 gpio_vtrip_sel[21]
port 806 nsew signal output
rlabel metal2 s 87600 953270 87656 953726 6 gpio_vtrip_sel[22]
port 807 nsew signal output
rlabel metal2 s 36200 953270 36256 953726 6 gpio_vtrip_sel[23]
port 808 nsew signal output
rlabel metal3 s -400 914192 60 914262 4 gpio_vtrip_sel[24]
port 809 nsew signal output
rlabel metal3 s -400 744392 60 744462 4 gpio_vtrip_sel[25]
port 810 nsew signal output
rlabel metal3 s -400 701192 60 701262 4 gpio_vtrip_sel[26]
port 811 nsew signal output
rlabel metal3 s -400 657992 60 658062 4 gpio_vtrip_sel[27]
port 812 nsew signal output
rlabel metal3 s -400 614792 60 614862 4 gpio_vtrip_sel[28]
port 813 nsew signal output
rlabel metal3 s -400 571592 60 571662 4 gpio_vtrip_sel[29]
port 814 nsew signal output
rlabel metal3 s 633266 161864 633726 161934 6 gpio_vtrip_sel[2]
port 815 nsew signal output
rlabel metal3 s -400 528392 60 528462 4 gpio_vtrip_sel[30]
port 816 nsew signal output
rlabel metal3 s -400 485192 60 485262 4 gpio_vtrip_sel[31]
port 817 nsew signal output
rlabel metal3 s -400 357592 60 357662 4 gpio_vtrip_sel[32]
port 818 nsew signal output
rlabel metal3 s -400 314392 60 314462 4 gpio_vtrip_sel[33]
port 819 nsew signal output
rlabel metal3 s -400 271192 60 271262 4 gpio_vtrip_sel[34]
port 820 nsew signal output
rlabel metal3 s -400 227992 60 228062 4 gpio_vtrip_sel[35]
port 821 nsew signal output
rlabel metal3 s -400 184792 60 184862 4 gpio_vtrip_sel[36]
port 822 nsew signal output
rlabel metal3 s -400 141592 60 141662 4 gpio_vtrip_sel[37]
port 823 nsew signal output
rlabel metal2 s 158070 -400 158126 56 8 gpio_vtrip_sel[38]
port 824 nsew signal output
rlabel metal2 s 266670 -400 266726 56 8 gpio_vtrip_sel[39]
port 825 nsew signal output
rlabel metal3 s 633266 207064 633726 207134 6 gpio_vtrip_sel[3]
port 826 nsew signal output
rlabel metal2 s 321470 -400 321526 56 8 gpio_vtrip_sel[40]
port 827 nsew signal output
rlabel metal2 s 376270 -400 376326 56 8 gpio_vtrip_sel[41]
port 828 nsew signal output
rlabel metal2 s 431070 -400 431126 56 8 gpio_vtrip_sel[42]
port 829 nsew signal output
rlabel metal2 s 485870 -400 485926 56 8 gpio_vtrip_sel[43]
port 830 nsew signal output
rlabel metal3 s 633266 252064 633726 252134 6 gpio_vtrip_sel[4]
port 831 nsew signal output
rlabel metal3 s 633266 297064 633726 297134 6 gpio_vtrip_sel[5]
port 832 nsew signal output
rlabel metal3 s 633266 342264 633726 342334 6 gpio_vtrip_sel[6]
port 833 nsew signal output
rlabel metal3 s 633266 519464 633726 519534 6 gpio_vtrip_sel[7]
port 834 nsew signal output
rlabel metal3 s 633266 564664 633726 564734 6 gpio_vtrip_sel[8]
port 835 nsew signal output
rlabel metal3 s 633266 609664 633726 609734 6 gpio_vtrip_sel[9]
port 836 nsew signal output
rlabel metal2 s 605082 -400 605134 56 8 mask_rev[0]
port 837 nsew signal input
rlabel metal2 s 607322 -400 607374 56 8 mask_rev[10]
port 838 nsew signal input
rlabel metal2 s 607546 -400 607598 56 8 mask_rev[11]
port 839 nsew signal input
rlabel metal2 s 607770 -400 607822 56 8 mask_rev[12]
port 840 nsew signal input
rlabel metal2 s 607994 -400 608046 56 8 mask_rev[13]
port 841 nsew signal input
rlabel metal2 s 608218 -400 608270 56 8 mask_rev[14]
port 842 nsew signal input
rlabel metal2 s 608442 -400 608494 56 8 mask_rev[15]
port 843 nsew signal input
rlabel metal2 s 608666 -400 608718 56 8 mask_rev[16]
port 844 nsew signal input
rlabel metal2 s 608890 -400 608942 56 8 mask_rev[17]
port 845 nsew signal input
rlabel metal2 s 609114 -400 609166 56 8 mask_rev[18]
port 846 nsew signal input
rlabel metal2 s 609338 -400 609390 56 8 mask_rev[19]
port 847 nsew signal input
rlabel metal2 s 605306 -400 605358 56 8 mask_rev[1]
port 848 nsew signal input
rlabel metal2 s 609562 -400 609614 56 8 mask_rev[20]
port 849 nsew signal input
rlabel metal2 s 609786 -400 609838 56 8 mask_rev[21]
port 850 nsew signal input
rlabel metal2 s 610010 -400 610062 56 8 mask_rev[22]
port 851 nsew signal input
rlabel metal2 s 610234 -400 610286 56 8 mask_rev[23]
port 852 nsew signal input
rlabel metal2 s 610458 -400 610510 56 8 mask_rev[24]
port 853 nsew signal input
rlabel metal2 s 610682 -400 610734 56 8 mask_rev[25]
port 854 nsew signal input
rlabel metal2 s 610906 -400 610958 56 8 mask_rev[26]
port 855 nsew signal input
rlabel metal2 s 611130 -400 611182 56 8 mask_rev[27]
port 856 nsew signal input
rlabel metal2 s 611354 -400 611406 56 8 mask_rev[28]
port 857 nsew signal input
rlabel metal2 s 611578 -400 611630 56 8 mask_rev[29]
port 858 nsew signal input
rlabel metal2 s 605530 -400 605582 56 8 mask_rev[2]
port 859 nsew signal input
rlabel metal2 s 611802 -400 611854 56 8 mask_rev[30]
port 860 nsew signal input
rlabel metal2 s 612026 -400 612078 56 8 mask_rev[31]
port 861 nsew signal input
rlabel metal2 s 605754 -400 605806 56 8 mask_rev[3]
port 862 nsew signal input
rlabel metal2 s 605978 -400 606030 56 8 mask_rev[4]
port 863 nsew signal input
rlabel metal2 s 606202 -400 606254 56 8 mask_rev[5]
port 864 nsew signal input
rlabel metal2 s 606426 -400 606478 56 8 mask_rev[6]
port 865 nsew signal input
rlabel metal2 s 606650 -400 606702 56 8 mask_rev[7]
port 866 nsew signal input
rlabel metal2 s 606874 -400 606926 56 8 mask_rev[8]
port 867 nsew signal input
rlabel metal2 s 607098 -400 607150 56 8 mask_rev[9]
port 868 nsew signal input
rlabel metal3 s -400 53372 60 53442 4 por_l
port 869 nsew signal input
rlabel metal3 s -400 53147 60 53217 4 porb_h
port 870 nsew signal input
rlabel metal3 s -400 53595 60 53665 4 porb_l
port 871 nsew signal input
rlabel metal2 s 99576 -400 99632 56 8 resetb_h
port 872 nsew signal input
rlabel metal2 s 110164 -400 110220 56 8 resetb_l
port 873 nsew signal input
rlabel metal3 s -400 25962 60 30762 4 vccd
port 874 nsew power input
rlabel metal3 s -400 36014 60 40804 4 vccd
port 874 nsew power input
rlabel metal3 s 633266 865522 633726 870312 6 vccd1
port 876 nsew power bidirectional
rlabel metal3 s 633266 875562 633726 880362 6 vccd1
port 876 nsew power bidirectional
rlabel metal3 s 633266 422810 633726 427472 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 4804 4960 8804 948128 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 4804 4960 628524 8960 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 4804 944128 628524 948128 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 624524 4960 628524 948128 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 11050 480 12330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 19050 480 20330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 27050 480 28330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 35050 480 36330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 43050 480 44330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 51050 480 52330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 59050 480 60330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 67050 480 68330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 75050 480 76330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 83050 480 84330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 91050 480 92330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 99050 480 100330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 107050 480 108330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 115050 480 116330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 123050 480 124330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 131050 480 132330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 139050 480 140330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 147050 480 148330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 155050 480 156330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 163050 480 164330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 171050 480 172330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 179050 480 180330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 187050 480 188330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 195050 480 196330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 203050 480 204330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 211050 480 212330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 219050 480 220330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 227050 480 228330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 235050 480 236330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 243050 480 244330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 251050 480 252330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 259050 480 260330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 267050 480 268330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 275050 480 276330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 283050 480 284330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 291050 480 292330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 299050 480 300330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 307050 480 308330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 315050 480 316330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 323050 480 324330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 331050 480 332330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 339050 480 340330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 347050 480 348330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 355050 480 356330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 363050 480 364330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 371050 480 372330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 379050 480 380330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 387050 480 388330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 395050 480 396330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 403050 480 404330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 411050 480 412330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 419050 480 420330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 427050 480 428330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 435050 480 436330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 443050 480 444330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 451050 480 452330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 459050 480 460330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 467050 480 468330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 475050 480 476330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 483050 480 484330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 491050 480 492330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 499050 480 500330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 507050 480 508330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 515050 480 516330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 523050 480 524330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 531050 480 532330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 539050 480 540330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 547050 480 548330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 555050 480 556330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 563050 480 564330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 571050 480 572330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 579050 480 580330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 587050 480 588330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 595050 480 596330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 603050 480 604330 57195 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 603050 372861 604330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 611050 480 612330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal4 s 619050 480 620330 952608 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 12086 633004 13366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 20086 633004 21366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 28086 633004 29366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 36086 633004 37366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 44086 633004 45366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 52086 633004 53366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 60086 633004 61366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 68086 633004 69366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 76086 633004 77366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 84086 633004 85366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 92086 633004 93366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 100086 633004 101366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 108086 633004 109366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 116086 633004 117366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 124086 633004 125366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 132086 633004 133366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 140086 633004 141366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 148086 633004 149366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 156086 633004 157366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 164086 633004 165366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 172086 633004 173366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 180086 633004 181366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 188086 633004 189366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 196086 633004 197366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 204086 633004 205366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 212086 633004 213366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 220086 633004 221366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 228086 633004 229366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 236086 633004 237366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 244086 633004 245366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 252086 633004 253366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 260086 633004 261366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 268086 633004 269366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 276086 633004 277366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 284086 633004 285366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 292086 633004 293366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 300086 633004 301366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 308086 633004 309366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 316086 633004 317366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 324086 633004 325366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 332086 633004 333366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 340086 633004 341366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 348086 633004 349366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 356086 633004 357366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 364086 633004 365366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 372086 633004 373366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 380086 633004 381366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 388086 633004 389366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 396086 633004 397366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 404086 633004 405366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 412086 633004 413366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 420086 633004 421366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 428086 633004 429366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 436086 633004 437366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 444086 633004 445366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 452086 633004 453366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 460086 633004 461366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 468086 633004 469366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 476086 633004 477366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 484086 633004 485366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 492086 633004 493366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 500086 633004 501366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 508086 633004 509366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 516086 633004 517366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 524086 633004 525366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 532086 633004 533366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 540086 633004 541366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 548086 633004 549366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 556086 633004 557366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 564086 633004 565366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 572086 633004 573366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 580086 633004 581366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 588086 633004 589366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 596086 633004 597366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 604086 633004 605366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 612086 633004 613366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 620086 633004 621366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 628086 633004 629366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 636086 633004 637366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 644086 633004 645366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 652086 633004 653366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 660086 633004 661366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 668086 633004 669366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 676086 633004 677366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 684086 633004 685366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 692086 633004 693366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 700086 633004 701366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 708086 633004 709366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 716086 633004 717366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 724086 633004 725366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 732086 633004 733366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 740086 633004 741366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 748086 633004 749366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 756086 633004 757366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 764086 633004 765366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 772086 633004 773366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 780086 633004 781366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 788086 633004 789366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 796086 633004 797366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 804086 633004 805366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 812086 633004 813366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 820086 633004 821366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 828086 633004 829366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 836086 633004 837366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 844086 633004 845366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 852086 633004 853366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 860086 633004 861366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 868086 633004 869366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 876086 633004 877366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 884086 633004 885366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 892086 633004 893366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 900086 633004 901366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 908086 633004 909366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 916086 633004 917366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 924086 633004 925366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 932086 633004 933366 6 vccd1
port 876 nsew power bidirectional
rlabel metal5 s 324 940086 633004 941366 6 vccd1
port 876 nsew power bidirectional
rlabel metal3 s -400 403862 60 408514 4 vccd2
port 880 nsew power input
rlabel metal3 s -400 869964 60 874764 4 vccd2
port 880 nsew power input
rlabel metal3 s -400 880014 60 884804 4 vccd2
port 880 nsew power input
rlabel metal3 s 580806 -400 585586 60 8 vdda
port 883 nsew power input
rlabel metal3 s 590784 -400 595564 60 8 vdda
port 883 nsew power input
rlabel metal3 s 633266 776406 633726 781186 6 vdda1
port 885 nsew power input
rlabel metal3 s 633266 461804 633726 466584 6 vdda1
port 885 nsew power input
rlabel metal3 s 633266 471784 633726 476564 6 vdda1
port 885 nsew power input
rlabel metal3 s 633266 786384 633726 791164 6 vdda1
port 885 nsew power input
rlabel metal3 s -400 450940 60 455720 4 vdda2
port 889 nsew power input
rlabel metal3 s -400 440962 60 445742 4 vdda2
port 889 nsew power input
rlabel metal3 s -400 78140 60 82920 4 vddio
port 891 nsew power input
rlabel metal3 s -400 837742 60 842522 4 vddio
port 891 nsew power input
rlabel metal3 s -400 68162 60 72942 4 vddio
port 891 nsew power input
rlabel metal3 s -400 827762 60 832542 4 vddio
port 891 nsew power input
rlabel metal3 s 46784 -400 51564 60 8 vssa
port 895 nsew ground input
rlabel metal3 s 36806 -400 41586 60 8 vssa
port 895 nsew ground input
rlabel metal3 s 543542 953266 548322 953726 6 vssa1
port 897 nsew ground input
rlabel metal3 s 633266 373606 633726 378386 6 vssa1
port 897 nsew ground input
rlabel metal3 s 533562 953266 538342 953726 6 vssa1
port 897 nsew ground input
rlabel metal3 s 633266 383584 633726 388364 6 vssa1
port 897 nsew ground input
rlabel metal3 s -400 795542 60 800322 4 vssa2
port 901 nsew ground input
rlabel metal3 s -400 785562 60 790342 4 vssa2
port 901 nsew ground input
rlabel metal3 s 209164 -400 213964 60 8 vssd
port 903 nsew ground input
rlabel metal3 s 199284 -400 203914 60 8 vssd
port 903 nsew ground input
rlabel metal3 s 633266 870610 633726 875272 6 vssd1
port 905 nsew ground bidirectional
rlabel metal3 s 633266 427762 633726 432562 6 vssd1
port 905 nsew ground bidirectional
rlabel metal3 s 633266 417722 633726 422512 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 324 480 4324 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 480 633004 4480 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 948608 633004 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 629004 480 633004 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 12970 480 14250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 20970 480 22250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 28970 480 30250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 36970 480 38250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 44970 480 46250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 52970 480 54250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 60970 480 62250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 68970 480 70250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 76970 480 78250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 84970 480 86250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 92970 480 94250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 100970 480 102250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 108970 480 110250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 116970 480 118250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 124970 480 126250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 132970 480 134250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 140970 480 142250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 148970 480 150250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 156970 480 158250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 164970 480 166250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 172970 480 174250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 180970 480 182250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 188970 480 190250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 196970 480 198250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 204970 480 206250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 212970 480 214250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 220970 480 222250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 228970 480 230250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 236970 480 238250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 244970 480 246250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 252970 480 254250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 260970 480 262250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 268970 480 270250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 276970 480 278250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 284970 480 286250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 292970 480 294250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 300970 480 302250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 308970 480 310250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 316970 480 318250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 324970 480 326250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 332970 480 334250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 340970 480 342250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 348970 480 350250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 356970 480 358250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 364970 480 366250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 372970 480 374250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 380970 480 382250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 388970 480 390250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 396970 480 398250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 404970 480 406250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 412970 480 414250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 420970 480 422250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 428970 480 430250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 436970 480 438250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 444970 480 446250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 452970 480 454250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 460970 480 462250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 468970 480 470250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 476970 480 478250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 484970 480 486250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 492970 480 494250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 500970 480 502250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 508970 480 510250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 516970 480 518250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 524970 480 526250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 532970 480 534250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 540970 480 542250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 548970 480 550250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 556970 480 558250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 564970 480 566250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 572970 480 574250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 580970 480 582250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 588970 480 590250 46988 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 588970 746596 590250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 596970 480 598250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 604970 480 606250 46988 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 604970 746596 606250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 612970 480 614250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal4 s 620970 480 622250 952608 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 14006 633004 15286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 22006 633004 23286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 30006 633004 31286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 38006 633004 39286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 46006 633004 47286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 54006 633004 55286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 62006 633004 63286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 70006 633004 71286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 78006 633004 79286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 86006 633004 87286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 94006 633004 95286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 102006 633004 103286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 110006 633004 111286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 118006 633004 119286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 126006 633004 127286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 134006 633004 135286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 142006 633004 143286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 150006 633004 151286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 158006 633004 159286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 166006 633004 167286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 174006 633004 175286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 182006 633004 183286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 190006 633004 191286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 198006 633004 199286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 206006 633004 207286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 214006 633004 215286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 222006 633004 223286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 230006 633004 231286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 238006 633004 239286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 246006 633004 247286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 254006 633004 255286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 262006 633004 263286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 270006 633004 271286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 278006 633004 279286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 286006 633004 287286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 294006 633004 295286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 302006 633004 303286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 310006 633004 311286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 318006 633004 319286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 326006 633004 327286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 334006 633004 335286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 342006 633004 343286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 350006 633004 351286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 358006 633004 359286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 366006 633004 367286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 374006 633004 375286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 382006 633004 383286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 390006 633004 391286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 398006 633004 399286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 406006 633004 407286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 414006 633004 415286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 422006 633004 423286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 430006 633004 431286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 438006 633004 439286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 446006 633004 447286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 454006 633004 455286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 462006 633004 463286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 470006 633004 471286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 478006 633004 479286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 486006 633004 487286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 494006 633004 495286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 502006 633004 503286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 510006 633004 511286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 518006 633004 519286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 526006 633004 527286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 534006 633004 535286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 542006 633004 543286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 550006 633004 551286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 558006 633004 559286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 566006 633004 567286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 574006 633004 575286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 582006 633004 583286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 590006 633004 591286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 598006 633004 599286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 606006 633004 607286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 614006 633004 615286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 622006 633004 623286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 630006 633004 631286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 638006 633004 639286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 646006 633004 647286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 654006 633004 655286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 662006 633004 663286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 670006 633004 671286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 678006 633004 679286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 686006 633004 687286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 694006 633004 695286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 702006 633004 703286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 710006 633004 711286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 718006 633004 719286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 726006 633004 727286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 734006 633004 735286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 742006 633004 743286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 750006 633004 751286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 758006 633004 759286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 766006 633004 767286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 774006 633004 775286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 782006 633004 783286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 790006 633004 791286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 798006 633004 799286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 806006 633004 807286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 814006 633004 815286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 822006 633004 823286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 830006 633004 831286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 838006 633004 839286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 846006 633004 847286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 854006 633004 855286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 862006 633004 863286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 870006 633004 871286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 878006 633004 879286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 886006 633004 887286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 894006 633004 895286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 902006 633004 903286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 910006 633004 911286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 918006 633004 919286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 926006 633004 927286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 934006 633004 935286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal5 s 324 942006 633004 943286 6 vssd1
port 905 nsew ground bidirectional
rlabel metal3 s -400 398762 60 403562 4 vssd2
port 909 nsew ground input
rlabel metal3 s -400 408814 60 413604 4 vssd2
port 909 nsew ground input
rlabel metal3 s -400 875054 60 879716 4 vssd2
port 909 nsew ground input
rlabel metal3 s 527006 -400 531786 60 8 vssio
port 912 nsew ground input
rlabel metal3 s 301342 953266 306122 953726 6 vssio
port 912 nsew ground input
rlabel metal3 s 536984 -400 541764 60 8 vssio
port 912 nsew ground input
rlabel metal3 s 291362 953266 296142 953726 6 vssio
port 912 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 633326 953326
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 31404248
string GDS_FILE /home/ghp7482/projects/LLM4Microwatt/openlane/openframe_project_wrapper/runs/25_10_21_14_31/results/signoff/openframe_project_wrapper.magic.gds
string GDS_START 10213156
<< end >>

